* File: Coin_bank.pex.sp
* Created: Wed Jan 17 12:36:35 2024
* Program "Calibre xRC"
* Version "v2021.3_35.19"
* 
.include "Coin_bank.pex.sp.pex"
.subckt COIN_BANK  VSS INIT3 INIT1 INIT0 STATE0 VDD STATE1 INIT2 POWER CLK STORE
+ MO2 MO0 MO3 MO1 M3 M1 M2 M0 S3 S2 S1 S0
* 
* S0	S0
* S1	S1
* S2	S2
* S3	S3
* M0	M0
* M2	M2
* M1	M1
* M3	M3
* MO1	MO1
* MO3	MO3
* MO0	MO0
* MO2	MO2
* STORE	STORE
* CLK	CLK
* POWER	POWER
* INIT2	INIT2
* STATE1	STATE1
* VDD	VDD
* STATE0	STATE0
* INIT0	INIT0
* INIT1	INIT1
* INIT3	INIT3
* VSS	VSS
mX0/M0 N_32_X0/M0_d N_STATE1_X0/M0_g N_VSS_X0/M0_s N_VSS_X0/M0_b N_18 L=1.8e-07
+ W=2.5e-06 AD=1.1625e-12 AS=2.325e-12 PD=9.3e-07 PS=4.36e-06
mX0/M1 N_VSS_X0/M1_d N_STATE1_X0/M1_g N_32_X0/M1_s N_VSS_X0/M0_b N_18 L=1.8e-07
+ W=2.5e-06 AD=1.95e-12 AS=1.1625e-12 PD=4.06e-06 PS=9.3e-07
mX0/M2 N_32_X0/M2_d N_STATE1_X0/M2_g N_VDD_X0/M2_s N_VDD_X0/M2_b P_18 L=1.8e-07
+ W=3e-06 AD=1.395e-12 AS=2.79e-12 PD=9.3e-07 PS=4.86e-06
mX0/M3 N_VDD_X0/M3_d N_STATE1_X0/M3_g N_32_X0/M3_s N_VDD_X0/M2_b P_18 L=1.8e-07
+ W=3e-06 AD=2.37e-12 AS=1.395e-12 PD=4.58e-06 PS=9.3e-07
mX1/M0 N_24_X1/M0_d N_STATE0_X1/M0_g N_VSS_X1/M0_s N_VSS_X0/M0_b N_18 L=1.8e-07
+ W=2.5e-06 AD=1.1625e-12 AS=2.325e-12 PD=9.3e-07 PS=4.36e-06
mX1/M1 N_VSS_X1/M1_d N_STATE0_X1/M1_g N_24_X1/M1_s N_VSS_X0/M0_b N_18 L=1.8e-07
+ W=2.5e-06 AD=1.95e-12 AS=1.1625e-12 PD=4.06e-06 PS=9.3e-07
mX1/M2 N_24_X1/M2_d N_STATE0_X1/M2_g N_VDD_X1/M2_s N_VDD_X1/M2_b P_18 L=1.8e-07
+ W=3e-06 AD=1.395e-12 AS=2.79e-12 PD=9.3e-07 PS=4.86e-06
mX1/M3 N_VDD_X1/M3_d N_STATE0_X1/M3_g N_24_X1/M3_s N_VDD_X1/M2_b P_18 L=1.8e-07
+ W=3e-06 AD=2.37e-12 AS=1.395e-12 PD=4.58e-06 PS=9.3e-07
mX2/M0 N_33_X2/M0_d N_STATE1_X2/M0_g N_VSS_X2/M0_s N_VSS_X0/M0_b N_18 L=1.8e-07
+ W=2.5e-06 AD=1.1625e-12 AS=2.325e-12 PD=9.3e-07 PS=4.36e-06
mX2/M1 N_VSS_X2/M1_d N_STATE1_X2/M1_g N_33_X2/M1_s N_VSS_X0/M0_b N_18 L=1.8e-07
+ W=2.5e-06 AD=1.95e-12 AS=1.1625e-12 PD=4.06e-06 PS=9.3e-07
mX2/M2 N_33_X2/M2_d N_STATE1_X2/M2_g N_VDD_X2/M2_s N_VDD_X2/M2_b P_18 L=1.8e-07
+ W=3e-06 AD=1.395e-12 AS=2.79e-12 PD=9.3e-07 PS=4.86e-06
mX2/M3 N_VDD_X2/M3_d N_STATE1_X2/M3_g N_33_X2/M3_s N_VDD_X2/M2_b P_18 L=1.8e-07
+ W=3e-06 AD=2.37e-12 AS=1.395e-12 PD=4.58e-06 PS=9.3e-07
mX3/M0 N_X3/9_X3/M0_d N_4_X3/M0_g N_VSS_X3/M0_s N_VSS_X0/M0_b N_18 L=1.8e-07
+ W=1.4e-06 AD=5.18e-13 AS=1.022e-12 PD=7.4e-07 PS=2.86e-06
mX3/M1 N_VSS_X3/M1_d N_INIT0_X3/M1_g N_X3/9_X3/M1_s N_VSS_X0/M0_b N_18 L=1.8e-07
+ W=1.4e-06 AD=9.24e-13 AS=5.18e-13 PD=2.72e-06 PS=7.4e-07
mX3/M2 N_X3/8_X3/M2_d N_VSS_X3/M2_g N_X3/9_X3/M2_s N_VSS_X0/M0_b N_18 L=1.8e-07
+ W=1.4e-06 AD=1.008e-12 AS=1.022e-12 PD=2.84e-06 PS=2.86e-06
mX3/M3 N_X3/17_X3/M3_d N_INIT0_X3/M3_g N_VSS_X3/M3_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=5.04e-13 AS=9.8e-13 PD=7.2e-07 PS=2.8e-06
mX3/M4 N_X3/8_X3/M4_d N_4_X3/M4_g N_X3/17_X3/M4_s N_VSS_X0/M0_b N_18 L=1.8e-07
+ W=1.4e-06 AD=9.94e-13 AS=5.04e-13 PD=2.82e-06 PS=7.2e-07
mX3/M5 N_X3/11_X3/M5_d N_4_X3/M5_g N_VSS_X3/M5_s N_VSS_X0/M0_b N_18 L=1.8e-07
+ W=1.4e-06 AD=4.83e-13 AS=1.12e-12 PD=6.9e-07 PS=3e-06
mX3/M6 N_VSS_X3/M6_d N_INIT0_X3/M6_g N_X3/11_X3/M6_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=5.6e-13 AS=4.83e-13 PD=8e-07 PS=6.9e-07
mX3/M7 N_X3/11_X3/M7_d N_VSS_X3/M7_g N_VSS_X3/M7_s N_VSS_X0/M0_b N_18 L=1.8e-07
+ W=1.4e-06 AD=1.022e-12 AS=5.6e-13 PD=2.86e-06 PS=8e-07
mX3/M8 N_X3/13_X3/M8_d N_X3/8_X3/M8_g N_X3/11_X3/M8_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=9.94e-13 AS=1.036e-12 PD=2.82e-06 PS=2.88e-06
mX3/M9 N_X3/18_X3/M9_d N_VSS_X3/M9_g N_VSS_X3/M9_s N_VSS_X0/M0_b N_18 L=1.8e-07
+ W=1.4e-06 AD=6.58e-13 AS=7.42e-13 PD=9.4e-07 PS=2.46e-06
mX3/M10 N_X3/19_X3/M10_d N_INIT0_X3/M10_g N_X3/18_X3/M10_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=6.44e-13 AS=6.58e-13 PD=9.2e-07 PS=9.4e-07
mX3/M11 N_X3/13_X3/M11_d N_4_X3/M11_g N_X3/19_X3/M11_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=8.82e-13 AS=6.44e-13 PD=2.66e-06 PS=9.2e-07
mX3/M12 N_X3/10_X3/M12_d N_4_X3/M12_g N_VDD_X3/M12_s N_VDD_X3/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=1.11e-12 AS=2.19e-12 PD=7.4e-07 PS=4.46e-06
mX3/M13 N_VDD_X3/M13_d N_INIT0_X3/M13_g N_X3/10_X3/M13_s N_VDD_X3/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=2.19e-12 AS=1.11e-12 PD=4.46e-06 PS=7.4e-07
mX3/M14 N_X3/8_X3/M14_d N_VSS_X3/M14_g N_X3/10_X3/M14_s N_VDD_X3/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=2.16e-12 AS=2.22e-12 PD=4.44e-06 PS=4.48e-06
mX3/M15 N_X3/14_X3/M15_d N_INIT0_X3/M15_g N_VDD_X3/M15_s N_VDD_X3/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=1.08e-12 AS=2.28e-12 PD=7.2e-07 PS=4.52e-06
mX3/M16 N_X3/8_X3/M16_d N_4_X3/M16_g N_X3/14_X3/M16_s N_VDD_X3/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=2.16e-12 AS=1.08e-12 PD=4.44e-06 PS=7.2e-07
mX3/M17 N_X3/12_X3/M17_d N_4_X3/M17_g N_VDD_X3/M17_s N_VDD_X3/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=1.035e-12 AS=2.43e-12 PD=6.9e-07 PS=4.62e-06
mX3/M18 N_VDD_X3/M18_d N_INIT0_X3/M18_g N_X3/12_X3/M18_s N_VDD_X3/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=1.2e-12 AS=1.035e-12 PD=8e-07 PS=6.9e-07
mX3/M19 N_X3/12_X3/M19_d N_VSS_X3/M19_g N_VDD_X3/M19_s N_VDD_X3/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=2.19e-12 AS=1.2e-12 PD=4.46e-06 PS=8e-07
mX3/M20 N_X3/13_X3/M20_d N_X3/8_X3/M20_g N_X3/12_X3/M20_s N_VDD_X3/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=2.07e-12 AS=2.31e-12 PD=4.38e-06 PS=4.54e-06
mX3/M21 N_X3/15_X3/M21_d N_VSS_X3/M21_g N_VDD_X3/M21_s N_VDD_X3/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=1.41e-12 AS=1.59e-12 PD=9.4e-07 PS=4.06e-06
mX3/M22 N_X3/16_X3/M22_d N_INIT0_X3/M22_g N_X3/15_X3/M22_s N_VDD_X3/X24/M2_b
+ P_18 L=1.8e-07 W=3e-06 AD=1.38e-12 AS=1.41e-12 PD=9.2e-07 PS=9.4e-07
mX3/M23 N_X3/13_X3/M23_d N_4_X3/M23_g N_X3/16_X3/M23_s N_VDD_X3/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=1.92e-12 AS=1.38e-12 PD=4.28e-06 PS=9.2e-07
mX3/X24/M0 N_15_X3/X24/M0_d N_X3/8_X3/X24/M0_g N_VSS_X3/X24/M0_s N_VSS_X0/M0_b
+ N_18 L=1.8e-07 W=2.5e-06 AD=1.1625e-12 AS=2.325e-12 PD=9.3e-07 PS=4.36e-06
mX3/X24/M1 N_VSS_X3/X24/M1_d N_X3/8_X3/X24/M1_g N_15_X3/X24/M1_s N_VSS_X0/M0_b
+ N_18 L=1.8e-07 W=2.5e-06 AD=1.95e-12 AS=1.1625e-12 PD=4.06e-06 PS=9.3e-07
mX3/X24/M2 N_15_X3/X24/M2_d N_X3/8_X3/X24/M2_g N_VDD_X3/X24/M2_s
+ N_VDD_X3/X24/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.395e-12 AS=2.79e-12 PD=9.3e-07
+ PS=4.86e-06
mX3/X24/M3 N_VDD_X3/X24/M3_d N_X3/8_X3/X24/M3_g N_15_X3/X24/M3_s
+ N_VDD_X3/X24/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.37e-12 AS=1.395e-12 PD=4.58e-06
+ PS=9.3e-07
mX3/X25/M0 N_5_X3/X25/M0_d N_X3/13_X3/X25/M0_g N_VSS_X3/X25/M0_s N_VSS_X0/M0_b
+ N_18 L=1.8e-07 W=2.5e-06 AD=1.1625e-12 AS=2.325e-12 PD=9.3e-07 PS=4.36e-06
mX3/X25/M1 N_VSS_X3/X25/M1_d N_X3/13_X3/X25/M1_g N_5_X3/X25/M1_s N_VSS_X0/M0_b
+ N_18 L=1.8e-07 W=2.5e-06 AD=1.95e-12 AS=1.1625e-12 PD=4.06e-06 PS=9.3e-07
mX3/X25/M2 N_5_X3/X25/M2_d N_X3/13_X3/X25/M2_g N_VDD_X3/X25/M2_s
+ N_VDD_X3/X24/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.395e-12 AS=2.79e-12 PD=9.3e-07
+ PS=4.86e-06
mX3/X25/M3 N_VDD_X3/X25/M3_d N_X3/13_X3/X25/M3_g N_5_X3/X25/M3_s
+ N_VDD_X3/X24/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.37e-12 AS=1.395e-12 PD=4.58e-06
+ PS=9.3e-07
mX4/M0 N_X4/9_X4/M0_d N_16_X4/M0_g N_VSS_X4/M0_s N_VSS_X0/M0_b N_18 L=1.8e-07
+ W=1.4e-06 AD=5.18e-13 AS=1.022e-12 PD=7.4e-07 PS=2.86e-06
mX4/M1 N_VSS_X4/M1_d N_INIT3_X4/M1_g N_X4/9_X4/M1_s N_VSS_X0/M0_b N_18 L=1.8e-07
+ W=1.4e-06 AD=9.24e-13 AS=5.18e-13 PD=2.72e-06 PS=7.4e-07
mX4/M2 N_X4/8_X4/M2_d N_18_X4/M2_g N_X4/9_X4/M2_s N_VSS_X0/M0_b N_18 L=1.8e-07
+ W=1.4e-06 AD=1.008e-12 AS=1.022e-12 PD=2.84e-06 PS=2.86e-06
mX4/M3 N_X4/17_X4/M3_d N_INIT3_X4/M3_g N_VSS_X4/M3_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=5.04e-13 AS=9.8e-13 PD=7.2e-07 PS=2.8e-06
mX4/M4 N_X4/8_X4/M4_d N_16_X4/M4_g N_X4/17_X4/M4_s N_VSS_X0/M0_b N_18 L=1.8e-07
+ W=1.4e-06 AD=9.94e-13 AS=5.04e-13 PD=2.82e-06 PS=7.2e-07
mX4/M5 N_X4/11_X4/M5_d N_16_X4/M5_g N_VSS_X4/M5_s N_VSS_X0/M0_b N_18 L=1.8e-07
+ W=1.4e-06 AD=4.83e-13 AS=1.12e-12 PD=6.9e-07 PS=3e-06
mX4/M6 N_VSS_X4/M6_d N_INIT3_X4/M6_g N_X4/11_X4/M6_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=5.6e-13 AS=4.83e-13 PD=8e-07 PS=6.9e-07
mX4/M7 N_X4/11_X4/M7_d N_18_X4/M7_g N_VSS_X4/M7_s N_VSS_X0/M0_b N_18 L=1.8e-07
+ W=1.4e-06 AD=1.022e-12 AS=5.6e-13 PD=2.86e-06 PS=8e-07
mX4/M8 N_X4/13_X4/M8_d N_X4/8_X4/M8_g N_X4/11_X4/M8_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=9.94e-13 AS=1.036e-12 PD=2.82e-06 PS=2.88e-06
mX4/M9 N_X4/18_X4/M9_d N_18_X4/M9_g N_VSS_X4/M9_s N_VSS_X0/M0_b N_18 L=1.8e-07
+ W=1.4e-06 AD=6.58e-13 AS=7.42e-13 PD=9.4e-07 PS=2.46e-06
mX4/M10 N_X4/19_X4/M10_d N_INIT3_X4/M10_g N_X4/18_X4/M10_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=6.44e-13 AS=6.58e-13 PD=9.2e-07 PS=9.4e-07
mX4/M11 N_X4/13_X4/M11_d N_16_X4/M11_g N_X4/19_X4/M11_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=8.82e-13 AS=6.44e-13 PD=2.66e-06 PS=9.2e-07
mX4/M12 N_X4/10_X4/M12_d N_16_X4/M12_g N_VDD_X4/M12_s N_VDD_X4/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=1.11e-12 AS=2.19e-12 PD=7.4e-07 PS=4.46e-06
mX4/M13 N_VDD_X4/M13_d N_INIT3_X4/M13_g N_X4/10_X4/M13_s N_VDD_X4/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=2.19e-12 AS=1.11e-12 PD=4.46e-06 PS=7.4e-07
mX4/M14 N_X4/8_X4/M14_d N_18_X4/M14_g N_X4/10_X4/M14_s N_VDD_X4/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=2.16e-12 AS=2.22e-12 PD=4.44e-06 PS=4.48e-06
mX4/M15 N_X4/14_X4/M15_d N_INIT3_X4/M15_g N_VDD_X4/M15_s N_VDD_X4/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=1.08e-12 AS=2.28e-12 PD=7.2e-07 PS=4.52e-06
mX4/M16 N_X4/8_X4/M16_d N_16_X4/M16_g N_X4/14_X4/M16_s N_VDD_X4/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=2.16e-12 AS=1.08e-12 PD=4.44e-06 PS=7.2e-07
mX4/M17 N_X4/12_X4/M17_d N_16_X4/M17_g N_VDD_X4/M17_s N_VDD_X4/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=1.035e-12 AS=2.43e-12 PD=6.9e-07 PS=4.62e-06
mX4/M18 N_VDD_X4/M18_d N_INIT3_X4/M18_g N_X4/12_X4/M18_s N_VDD_X4/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=1.2e-12 AS=1.035e-12 PD=8e-07 PS=6.9e-07
mX4/M19 N_X4/12_X4/M19_d N_18_X4/M19_g N_VDD_X4/M19_s N_VDD_X4/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=2.19e-12 AS=1.2e-12 PD=4.46e-06 PS=8e-07
mX4/M20 N_X4/13_X4/M20_d N_X4/8_X4/M20_g N_X4/12_X4/M20_s N_VDD_X4/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=2.07e-12 AS=2.31e-12 PD=4.38e-06 PS=4.54e-06
mX4/M21 N_X4/15_X4/M21_d N_18_X4/M21_g N_VDD_X4/M21_s N_VDD_X4/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=1.41e-12 AS=1.59e-12 PD=9.4e-07 PS=4.06e-06
mX4/M22 N_X4/16_X4/M22_d N_INIT3_X4/M22_g N_X4/15_X4/M22_s N_VDD_X4/X24/M2_b
+ P_18 L=1.8e-07 W=3e-06 AD=1.38e-12 AS=1.41e-12 PD=9.2e-07 PS=9.4e-07
mX4/M23 N_X4/13_X4/M23_d N_16_X4/M23_g N_X4/16_X4/M23_s N_VDD_X4/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=1.92e-12 AS=1.38e-12 PD=4.28e-06 PS=9.2e-07
mX4/X24/M0 N_34_X4/X24/M0_d N_X4/8_X4/X24/M0_g N_VSS_X4/X24/M0_s N_VSS_X0/M0_b
+ N_18 L=1.8e-07 W=2.5e-06 AD=1.1625e-12 AS=2.325e-12 PD=9.3e-07 PS=4.36e-06
mX4/X24/M1 N_VSS_X4/X24/M1_d N_X4/8_X4/X24/M1_g N_34_X4/X24/M1_s N_VSS_X0/M0_b
+ N_18 L=1.8e-07 W=2.5e-06 AD=1.95e-12 AS=1.1625e-12 PD=4.06e-06 PS=9.3e-07
mX4/X24/M2 N_34_X4/X24/M2_d N_X4/8_X4/X24/M2_g N_VDD_X4/X24/M2_s
+ N_VDD_X4/X24/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.395e-12 AS=2.79e-12 PD=9.3e-07
+ PS=4.86e-06
mX4/X24/M3 N_VDD_X4/X24/M3_d N_X4/8_X4/X24/M3_g N_34_X4/X24/M3_s
+ N_VDD_X4/X24/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.37e-12 AS=1.395e-12 PD=4.58e-06
+ PS=9.3e-07
mX4/X25/M0 N_14_X4/X25/M0_d N_X4/13_X4/X25/M0_g N_VSS_X4/X25/M0_s N_VSS_X0/M0_b
+ N_18 L=1.8e-07 W=2.5e-06 AD=1.1625e-12 AS=2.325e-12 PD=9.3e-07 PS=4.36e-06
mX4/X25/M1 N_VSS_X4/X25/M1_d N_X4/13_X4/X25/M1_g N_14_X4/X25/M1_s N_VSS_X0/M0_b
+ N_18 L=1.8e-07 W=2.5e-06 AD=1.95e-12 AS=1.1625e-12 PD=4.06e-06 PS=9.3e-07
mX4/X25/M2 N_14_X4/X25/M2_d N_X4/13_X4/X25/M2_g N_VDD_X4/X25/M2_s
+ N_VDD_X4/X24/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.395e-12 AS=2.79e-12 PD=9.3e-07
+ PS=4.86e-06
mX4/X25/M3 N_VDD_X4/X25/M3_d N_X4/13_X4/X25/M3_g N_14_X4/X25/M3_s
+ N_VDD_X4/X24/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.37e-12 AS=1.395e-12 PD=4.58e-06
+ PS=9.3e-07
mX5/M0 N_X5/9_X5/M0_d N_10_X5/M0_g N_VSS_X5/M0_s N_VSS_X0/M0_b N_18 L=1.8e-07
+ W=1.4e-06 AD=5.18e-13 AS=1.022e-12 PD=7.4e-07 PS=2.86e-06
mX5/M1 N_VSS_X5/M1_d N_INIT1_X5/M1_g N_X5/9_X5/M1_s N_VSS_X0/M0_b N_18 L=1.8e-07
+ W=1.4e-06 AD=9.24e-13 AS=5.18e-13 PD=2.72e-06 PS=7.4e-07
mX5/M2 N_X5/8_X5/M2_d N_15_X5/M2_g N_X5/9_X5/M2_s N_VSS_X0/M0_b N_18 L=1.8e-07
+ W=1.4e-06 AD=1.008e-12 AS=1.022e-12 PD=2.84e-06 PS=2.86e-06
mX5/M3 N_X5/17_X5/M3_d N_INIT1_X5/M3_g N_VSS_X5/M3_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=5.04e-13 AS=9.8e-13 PD=7.2e-07 PS=2.8e-06
mX5/M4 N_X5/8_X5/M4_d N_10_X5/M4_g N_X5/17_X5/M4_s N_VSS_X0/M0_b N_18 L=1.8e-07
+ W=1.4e-06 AD=9.94e-13 AS=5.04e-13 PD=2.82e-06 PS=7.2e-07
mX5/M5 N_X5/11_X5/M5_d N_10_X5/M5_g N_VSS_X5/M5_s N_VSS_X0/M0_b N_18 L=1.8e-07
+ W=1.4e-06 AD=4.83e-13 AS=1.12e-12 PD=6.9e-07 PS=3e-06
mX5/M6 N_VSS_X5/M6_d N_INIT1_X5/M6_g N_X5/11_X5/M6_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=5.6e-13 AS=4.83e-13 PD=8e-07 PS=6.9e-07
mX5/M7 N_X5/11_X5/M7_d N_15_X5/M7_g N_VSS_X5/M7_s N_VSS_X0/M0_b N_18 L=1.8e-07
+ W=1.4e-06 AD=1.022e-12 AS=5.6e-13 PD=2.86e-06 PS=8e-07
mX5/M8 N_X5/13_X5/M8_d N_X5/8_X5/M8_g N_X5/11_X5/M8_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=9.94e-13 AS=1.036e-12 PD=2.82e-06 PS=2.88e-06
mX5/M9 N_X5/18_X5/M9_d N_15_X5/M9_g N_VSS_X5/M9_s N_VSS_X0/M0_b N_18 L=1.8e-07
+ W=1.4e-06 AD=6.58e-13 AS=7.42e-13 PD=9.4e-07 PS=2.46e-06
mX5/M10 N_X5/19_X5/M10_d N_INIT1_X5/M10_g N_X5/18_X5/M10_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=6.44e-13 AS=6.58e-13 PD=9.2e-07 PS=9.4e-07
mX5/M11 N_X5/13_X5/M11_d N_10_X5/M11_g N_X5/19_X5/M11_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=8.82e-13 AS=6.44e-13 PD=2.66e-06 PS=9.2e-07
mX5/M12 N_X5/10_X5/M12_d N_10_X5/M12_g N_VDD_X5/M12_s N_VDD_X3/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=1.11e-12 AS=2.19e-12 PD=7.4e-07 PS=4.46e-06
mX5/M13 N_VDD_X5/M13_d N_INIT1_X5/M13_g N_X5/10_X5/M13_s N_VDD_X3/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=2.19e-12 AS=1.11e-12 PD=4.46e-06 PS=7.4e-07
mX5/M14 N_X5/8_X5/M14_d N_15_X5/M14_g N_X5/10_X5/M14_s N_VDD_X3/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=2.16e-12 AS=2.22e-12 PD=4.44e-06 PS=4.48e-06
mX5/M15 N_X5/14_X5/M15_d N_INIT1_X5/M15_g N_VDD_X5/M15_s N_VDD_X3/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=1.08e-12 AS=2.28e-12 PD=7.2e-07 PS=4.52e-06
mX5/M16 N_X5/8_X5/M16_d N_10_X5/M16_g N_X5/14_X5/M16_s N_VDD_X3/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=2.16e-12 AS=1.08e-12 PD=4.44e-06 PS=7.2e-07
mX5/M17 N_X5/12_X5/M17_d N_10_X5/M17_g N_VDD_X5/M17_s N_VDD_X3/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=1.035e-12 AS=2.43e-12 PD=6.9e-07 PS=4.62e-06
mX5/M18 N_VDD_X5/M18_d N_INIT1_X5/M18_g N_X5/12_X5/M18_s N_VDD_X3/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=1.2e-12 AS=1.035e-12 PD=8e-07 PS=6.9e-07
mX5/M19 N_X5/12_X5/M19_d N_15_X5/M19_g N_VDD_X5/M19_s N_VDD_X3/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=2.19e-12 AS=1.2e-12 PD=4.46e-06 PS=8e-07
mX5/M20 N_X5/13_X5/M20_d N_X5/8_X5/M20_g N_X5/12_X5/M20_s N_VDD_X3/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=2.07e-12 AS=2.31e-12 PD=4.38e-06 PS=4.54e-06
mX5/M21 N_X5/15_X5/M21_d N_15_X5/M21_g N_VDD_X5/M21_s N_VDD_X3/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=1.41e-12 AS=1.59e-12 PD=9.4e-07 PS=4.06e-06
mX5/M22 N_X5/16_X5/M22_d N_INIT1_X5/M22_g N_X5/15_X5/M22_s N_VDD_X3/X24/M2_b
+ P_18 L=1.8e-07 W=3e-06 AD=1.38e-12 AS=1.41e-12 PD=9.2e-07 PS=9.4e-07
mX5/M23 N_X5/13_X5/M23_d N_10_X5/M23_g N_X5/16_X5/M23_s N_VDD_X3/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=1.92e-12 AS=1.38e-12 PD=4.28e-06 PS=9.2e-07
mX5/X24/M0 N_17_X5/X24/M0_d N_X5/8_X5/X24/M0_g N_VSS_X5/X24/M0_s N_VSS_X0/M0_b
+ N_18 L=1.8e-07 W=2.5e-06 AD=1.1625e-12 AS=2.325e-12 PD=9.3e-07 PS=4.36e-06
mX5/X24/M1 N_VSS_X5/X24/M1_d N_X5/8_X5/X24/M1_g N_17_X5/X24/M1_s N_VSS_X0/M0_b
+ N_18 L=1.8e-07 W=2.5e-06 AD=1.95e-12 AS=1.1625e-12 PD=4.06e-06 PS=9.3e-07
mX5/X24/M2 N_17_X5/X24/M2_d N_X5/8_X5/X24/M2_g N_VDD_X5/X24/M2_s
+ N_VDD_X3/X24/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.395e-12 AS=2.79e-12 PD=9.3e-07
+ PS=4.86e-06
mX5/X24/M3 N_VDD_X5/X24/M3_d N_X5/8_X5/X24/M3_g N_17_X5/X24/M3_s
+ N_VDD_X3/X24/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.37e-12 AS=1.395e-12 PD=4.58e-06
+ PS=9.3e-07
mX5/X25/M0 N_13_X5/X25/M0_d N_X5/13_X5/X25/M0_g N_VSS_X5/X25/M0_s N_VSS_X0/M0_b
+ N_18 L=1.8e-07 W=2.5e-06 AD=1.1625e-12 AS=2.325e-12 PD=9.3e-07 PS=4.36e-06
mX5/X25/M1 N_VSS_X5/X25/M1_d N_X5/13_X5/X25/M1_g N_13_X5/X25/M1_s N_VSS_X0/M0_b
+ N_18 L=1.8e-07 W=2.5e-06 AD=1.95e-12 AS=1.1625e-12 PD=4.06e-06 PS=9.3e-07
mX5/X25/M2 N_13_X5/X25/M2_d N_X5/13_X5/X25/M2_g N_VDD_X5/X25/M2_s
+ N_VDD_X3/X24/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.395e-12 AS=2.79e-12 PD=9.3e-07
+ PS=4.86e-06
mX5/X25/M3 N_VDD_X5/X25/M3_d N_X5/13_X5/X25/M3_g N_13_X5/X25/M3_s
+ N_VDD_X3/X24/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.37e-12 AS=1.395e-12 PD=4.58e-06
+ PS=9.3e-07
mX6/M0 N_X6/9_X6/M0_d N_3_X6/M0_g N_VSS_X6/M0_s N_VSS_X0/M0_b N_18 L=1.8e-07
+ W=1.4e-06 AD=5.18e-13 AS=1.022e-12 PD=7.4e-07 PS=2.86e-06
mX6/M1 N_VSS_X6/M1_d N_INIT2_X6/M1_g N_X6/9_X6/M1_s N_VSS_X0/M0_b N_18 L=1.8e-07
+ W=1.4e-06 AD=9.24e-13 AS=5.18e-13 PD=2.72e-06 PS=7.4e-07
mX6/M2 N_X6/8_X6/M2_d N_17_X6/M2_g N_X6/9_X6/M2_s N_VSS_X0/M0_b N_18 L=1.8e-07
+ W=1.4e-06 AD=1.008e-12 AS=1.022e-12 PD=2.84e-06 PS=2.86e-06
mX6/M3 N_X6/17_X6/M3_d N_INIT2_X6/M3_g N_VSS_X6/M3_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=5.04e-13 AS=9.8e-13 PD=7.2e-07 PS=2.8e-06
mX6/M4 N_X6/8_X6/M4_d N_3_X6/M4_g N_X6/17_X6/M4_s N_VSS_X0/M0_b N_18 L=1.8e-07
+ W=1.4e-06 AD=9.94e-13 AS=5.04e-13 PD=2.82e-06 PS=7.2e-07
mX6/M5 N_X6/11_X6/M5_d N_3_X6/M5_g N_VSS_X6/M5_s N_VSS_X0/M0_b N_18 L=1.8e-07
+ W=1.4e-06 AD=4.83e-13 AS=1.12e-12 PD=6.9e-07 PS=3e-06
mX6/M6 N_VSS_X6/M6_d N_INIT2_X6/M6_g N_X6/11_X6/M6_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=5.6e-13 AS=4.83e-13 PD=8e-07 PS=6.9e-07
mX6/M7 N_X6/11_X6/M7_d N_17_X6/M7_g N_VSS_X6/M7_s N_VSS_X0/M0_b N_18 L=1.8e-07
+ W=1.4e-06 AD=1.022e-12 AS=5.6e-13 PD=2.86e-06 PS=8e-07
mX6/M8 N_X6/13_X6/M8_d N_X6/8_X6/M8_g N_X6/11_X6/M8_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=9.94e-13 AS=1.036e-12 PD=2.82e-06 PS=2.88e-06
mX6/M9 N_X6/18_X6/M9_d N_17_X6/M9_g N_VSS_X6/M9_s N_VSS_X0/M0_b N_18 L=1.8e-07
+ W=1.4e-06 AD=6.58e-13 AS=7.42e-13 PD=9.4e-07 PS=2.46e-06
mX6/M10 N_X6/19_X6/M10_d N_INIT2_X6/M10_g N_X6/18_X6/M10_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=6.44e-13 AS=6.58e-13 PD=9.2e-07 PS=9.4e-07
mX6/M11 N_X6/13_X6/M11_d N_3_X6/M11_g N_X6/19_X6/M11_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=8.82e-13 AS=6.44e-13 PD=2.66e-06 PS=9.2e-07
mX6/M12 N_X6/10_X6/M12_d N_3_X6/M12_g N_VDD_X6/M12_s N_VDD_X4/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=1.11e-12 AS=2.19e-12 PD=7.4e-07 PS=4.46e-06
mX6/M13 N_VDD_X6/M13_d N_INIT2_X6/M13_g N_X6/10_X6/M13_s N_VDD_X4/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=2.19e-12 AS=1.11e-12 PD=4.46e-06 PS=7.4e-07
mX6/M14 N_X6/8_X6/M14_d N_17_X6/M14_g N_X6/10_X6/M14_s N_VDD_X4/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=2.16e-12 AS=2.22e-12 PD=4.44e-06 PS=4.48e-06
mX6/M15 N_X6/14_X6/M15_d N_INIT2_X6/M15_g N_VDD_X6/M15_s N_VDD_X4/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=1.08e-12 AS=2.28e-12 PD=7.2e-07 PS=4.52e-06
mX6/M16 N_X6/8_X6/M16_d N_3_X6/M16_g N_X6/14_X6/M16_s N_VDD_X4/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=2.16e-12 AS=1.08e-12 PD=4.44e-06 PS=7.2e-07
mX6/M17 N_X6/12_X6/M17_d N_3_X6/M17_g N_VDD_X6/M17_s N_VDD_X4/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=1.035e-12 AS=2.43e-12 PD=6.9e-07 PS=4.62e-06
mX6/M18 N_VDD_X6/M18_d N_INIT2_X6/M18_g N_X6/12_X6/M18_s N_VDD_X4/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=1.2e-12 AS=1.035e-12 PD=8e-07 PS=6.9e-07
mX6/M19 N_X6/12_X6/M19_d N_17_X6/M19_g N_VDD_X6/M19_s N_VDD_X4/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=2.19e-12 AS=1.2e-12 PD=4.46e-06 PS=8e-07
mX6/M20 N_X6/13_X6/M20_d N_X6/8_X6/M20_g N_X6/12_X6/M20_s N_VDD_X4/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=2.07e-12 AS=2.31e-12 PD=4.38e-06 PS=4.54e-06
mX6/M21 N_X6/15_X6/M21_d N_17_X6/M21_g N_VDD_X6/M21_s N_VDD_X4/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=1.41e-12 AS=1.59e-12 PD=9.4e-07 PS=4.06e-06
mX6/M22 N_X6/16_X6/M22_d N_INIT2_X6/M22_g N_X6/15_X6/M22_s N_VDD_X4/X24/M2_b
+ P_18 L=1.8e-07 W=3e-06 AD=1.38e-12 AS=1.41e-12 PD=9.2e-07 PS=9.4e-07
mX6/M23 N_X6/13_X6/M23_d N_3_X6/M23_g N_X6/16_X6/M23_s N_VDD_X4/X24/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=1.92e-12 AS=1.38e-12 PD=4.28e-06 PS=9.2e-07
mX6/X24/M0 N_18_X6/X24/M0_d N_X6/8_X6/X24/M0_g N_VSS_X6/X24/M0_s N_VSS_X0/M0_b
+ N_18 L=1.8e-07 W=2.5e-06 AD=1.1625e-12 AS=2.325e-12 PD=9.3e-07 PS=4.36e-06
mX6/X24/M1 N_VSS_X6/X24/M1_d N_X6/8_X6/X24/M1_g N_18_X6/X24/M1_s N_VSS_X0/M0_b
+ N_18 L=1.8e-07 W=2.5e-06 AD=1.95e-12 AS=1.1625e-12 PD=4.06e-06 PS=9.3e-07
mX6/X24/M2 N_18_X6/X24/M2_d N_X6/8_X6/X24/M2_g N_VDD_X6/X24/M2_s
+ N_VDD_X4/X24/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.395e-12 AS=2.79e-12 PD=9.3e-07
+ PS=4.86e-06
mX6/X24/M3 N_VDD_X6/X24/M3_d N_X6/8_X6/X24/M3_g N_18_X6/X24/M3_s
+ N_VDD_X4/X24/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.37e-12 AS=1.395e-12 PD=4.58e-06
+ PS=9.3e-07
mX6/X25/M0 N_27_X6/X25/M0_d N_X6/13_X6/X25/M0_g N_VSS_X6/X25/M0_s N_VSS_X0/M0_b
+ N_18 L=1.8e-07 W=2.5e-06 AD=1.1625e-12 AS=2.325e-12 PD=9.3e-07 PS=4.36e-06
mX6/X25/M1 N_VSS_X6/X25/M1_d N_X6/13_X6/X25/M1_g N_27_X6/X25/M1_s N_VSS_X0/M0_b
+ N_18 L=1.8e-07 W=2.5e-06 AD=1.95e-12 AS=1.1625e-12 PD=4.06e-06 PS=9.3e-07
mX6/X25/M2 N_27_X6/X25/M2_d N_X6/13_X6/X25/M2_g N_VDD_X6/X25/M2_s
+ N_VDD_X4/X24/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.395e-12 AS=2.79e-12 PD=9.3e-07
+ PS=4.86e-06
mX6/X25/M3 N_VDD_X6/X25/M3_d N_X6/13_X6/X25/M3_g N_27_X6/X25/M3_s
+ N_VDD_X4/X24/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.37e-12 AS=1.395e-12 PD=4.58e-06
+ PS=9.3e-07
mX7/X0/X0/M0 N_X7/X0/7_X7/X0/X0/M0_d N_STATE0_X7/X0/X0/M0_g N_VSS_X7/X0/X0/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.1625e-12 AS=2.325e-12 PD=9.3e-07
+ PS=4.36e-06
mX7/X0/X0/M1 N_VSS_X7/X0/X0/M1_d N_STATE0_X7/X0/X0/M1_g N_X7/X0/7_X7/X0/X0/M1_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.95e-12 AS=1.1625e-12 PD=4.06e-06
+ PS=9.3e-07
mX7/X0/X0/M2 N_X7/X0/7_X7/X0/X0/M2_d N_STATE0_X7/X0/X0/M2_g N_VDD_X7/X0/X0/M2_s
+ N_VDD_X7/X0/X0/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.395e-12 AS=2.79e-12 PD=9.3e-07
+ PS=4.86e-06
mX7/X0/X0/M3 N_VDD_X7/X0/X0/M3_d N_STATE0_X7/X0/X0/M3_g N_X7/X0/7_X7/X0/X0/M3_s
+ N_VDD_X7/X0/X0/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.37e-12 AS=1.395e-12
+ PD=4.58e-06 PS=9.3e-07
mX7/X0/X1/M0 N_X7/8_X7/X0/X1/M0_d N_STATE0_X7/X0/X1/M0_g N_INIT2_X7/X0/X1/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.316e-12 AS=1.288e-12 PD=3.28e-06
+ PS=3.24e-06
mX7/X0/X1/M1 N_X7/8_X7/X0/X1/M1_d N_X7/X0/7_X7/X0/X1/M1_g N_INIT2_X7/X0/X1/M1_s
+ N_VDD_X7/X0/X0/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.88e-12 AS=2.7e-12 PD=4.92e-06
+ PS=4.8e-06
mX7/X0/X2/M0 N_X7/8_X7/X0/X2/M0_d N_X7/X0/7_X7/X0/X2/M0_g N_3_X7/X0/X2/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.316e-12 AS=1.288e-12 PD=3.28e-06
+ PS=3.24e-06
mX7/X0/X2/M1 N_X7/8_X7/X0/X2/M1_d N_STATE0_X7/X0/X2/M1_g N_3_X7/X0/X2/M1_s
+ N_VDD_X7/X0/X0/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.88e-12 AS=2.7e-12 PD=4.92e-06
+ PS=4.8e-06
mX7/X1/X0/M0 N_X7/X1/7_X7/X1/X0/M0_d N_STATE1_X7/X1/X0/M0_g N_VSS_X7/X1/X0/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.1625e-12 AS=2.325e-12 PD=9.3e-07
+ PS=4.36e-06
mX7/X1/X0/M1 N_VSS_X7/X1/X0/M1_d N_STATE1_X7/X1/X0/M1_g N_X7/X1/7_X7/X1/X0/M1_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.95e-12 AS=1.1625e-12 PD=4.06e-06
+ PS=9.3e-07
mX7/X1/X0/M2 N_X7/X1/7_X7/X1/X0/M2_d N_STATE1_X7/X1/X0/M2_g N_VDD_X7/X1/X0/M2_s
+ N_VDD_X7/X0/X0/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.395e-12 AS=2.79e-12 PD=9.3e-07
+ PS=4.86e-06
mX7/X1/X0/M3 N_VDD_X7/X1/X0/M3_d N_STATE1_X7/X1/X0/M3_g N_X7/X1/7_X7/X1/X0/M3_s
+ N_VDD_X7/X0/X0/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.37e-12 AS=1.395e-12
+ PD=4.58e-06 PS=9.3e-07
mX7/X1/X1/M0 N_MO2_X7/X1/X1/M0_d N_STATE1_X7/X1/X1/M0_g N_X7/8_X7/X1/X1/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.316e-12 AS=1.288e-12 PD=3.28e-06
+ PS=3.24e-06
mX7/X1/X1/M1 N_MO2_X7/X1/X1/M1_d N_X7/X1/7_X7/X1/X1/M1_g N_X7/8_X7/X1/X1/M1_s
+ N_VDD_X7/X0/X0/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.88e-12 AS=2.7e-12 PD=4.92e-06
+ PS=4.8e-06
mX7/X1/X2/M0 N_MO2_X7/X1/X2/M0_d N_X7/X1/7_X7/X1/X2/M0_g N_VSS_X7/X1/X2/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.316e-12 AS=1.288e-12 PD=3.28e-06
+ PS=3.24e-06
mX7/X1/X2/M1 N_MO2_X7/X1/X2/M1_d N_STATE1_X7/X1/X2/M1_g N_VSS_X7/X1/X2/M1_s
+ N_VDD_X7/X0/X0/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.88e-12 AS=2.7e-12 PD=4.92e-06
+ PS=4.8e-06
mX8/X0/X0/M0 N_X8/X0/7_X8/X0/X0/M0_d N_STATE0_X8/X0/X0/M0_g N_VSS_X8/X0/X0/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.1625e-12 AS=2.325e-12 PD=9.3e-07
+ PS=4.36e-06
mX8/X0/X0/M1 N_VSS_X8/X0/X0/M1_d N_STATE0_X8/X0/X0/M1_g N_X8/X0/7_X8/X0/X0/M1_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.95e-12 AS=1.1625e-12 PD=4.06e-06
+ PS=9.3e-07
mX8/X0/X0/M2 N_X8/X0/7_X8/X0/X0/M2_d N_STATE0_X8/X0/X0/M2_g N_VDD_X8/X0/X0/M2_s
+ N_VDD_X2/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.395e-12 AS=2.79e-12 PD=9.3e-07
+ PS=4.86e-06
mX8/X0/X0/M3 N_VDD_X8/X0/X0/M3_d N_STATE0_X8/X0/X0/M3_g N_X8/X0/7_X8/X0/X0/M3_s
+ N_VDD_X2/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.37e-12 AS=1.395e-12 PD=4.58e-06
+ PS=9.3e-07
mX8/X0/X1/M0 N_X8/8_X8/X0/X1/M0_d N_STATE0_X8/X0/X1/M0_g N_INIT0_X8/X0/X1/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.316e-12 AS=1.288e-12 PD=3.28e-06
+ PS=3.24e-06
mX8/X0/X1/M1 N_X8/8_X8/X0/X1/M1_d N_X8/X0/7_X8/X0/X1/M1_g N_INIT0_X8/X0/X1/M1_s
+ N_VDD_X2/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.88e-12 AS=2.7e-12 PD=4.92e-06
+ PS=4.8e-06
mX8/X0/X2/M0 N_X8/8_X8/X0/X2/M0_d N_X8/X0/7_X8/X0/X2/M0_g N_4_X8/X0/X2/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.316e-12 AS=1.288e-12 PD=3.28e-06
+ PS=3.24e-06
mX8/X0/X2/M1 N_X8/8_X8/X0/X2/M1_d N_STATE0_X8/X0/X2/M1_g N_4_X8/X0/X2/M1_s
+ N_VDD_X2/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.88e-12 AS=2.7e-12 PD=4.92e-06
+ PS=4.8e-06
mX8/X1/X0/M0 N_X8/X1/7_X8/X1/X0/M0_d N_STATE1_X8/X1/X0/M0_g N_VSS_X8/X1/X0/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.1625e-12 AS=2.325e-12 PD=9.3e-07
+ PS=4.36e-06
mX8/X1/X0/M1 N_VSS_X8/X1/X0/M1_d N_STATE1_X8/X1/X0/M1_g N_X8/X1/7_X8/X1/X0/M1_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.95e-12 AS=1.1625e-12 PD=4.06e-06
+ PS=9.3e-07
mX8/X1/X0/M2 N_X8/X1/7_X8/X1/X0/M2_d N_STATE1_X8/X1/X0/M2_g N_VDD_X8/X1/X0/M2_s
+ N_VDD_X2/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.395e-12 AS=2.79e-12 PD=9.3e-07
+ PS=4.86e-06
mX8/X1/X0/M3 N_VDD_X8/X1/X0/M3_d N_STATE1_X8/X1/X0/M3_g N_X8/X1/7_X8/X1/X0/M3_s
+ N_VDD_X2/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.37e-12 AS=1.395e-12 PD=4.58e-06
+ PS=9.3e-07
mX8/X1/X1/M0 N_MO0_X8/X1/X1/M0_d N_STATE1_X8/X1/X1/M0_g N_X8/8_X8/X1/X1/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.316e-12 AS=1.288e-12 PD=3.28e-06
+ PS=3.24e-06
mX8/X1/X1/M1 N_MO0_X8/X1/X1/M1_d N_X8/X1/7_X8/X1/X1/M1_g N_X8/8_X8/X1/X1/M1_s
+ N_VDD_X2/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.88e-12 AS=2.7e-12 PD=4.92e-06
+ PS=4.8e-06
mX8/X1/X2/M0 N_MO0_X8/X1/X2/M0_d N_X8/X1/7_X8/X1/X2/M0_g N_VSS_X8/X1/X2/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.316e-12 AS=1.288e-12 PD=3.28e-06
+ PS=3.24e-06
mX8/X1/X2/M1 N_MO0_X8/X1/X2/M1_d N_STATE1_X8/X1/X2/M1_g N_VSS_X8/X1/X2/M1_s
+ N_VDD_X2/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.88e-12 AS=2.7e-12 PD=4.92e-06
+ PS=4.8e-06
mX9/X0/X0/M0 N_X9/X0/7_X9/X0/X0/M0_d N_STATE0_X9/X0/X0/M0_g N_VSS_X9/X0/X0/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.1625e-12 AS=2.325e-12 PD=9.3e-07
+ PS=4.36e-06
mX9/X0/X0/M1 N_VSS_X9/X0/X0/M1_d N_STATE0_X9/X0/X0/M1_g N_X9/X0/7_X9/X0/X0/M1_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.95e-12 AS=1.1625e-12 PD=4.06e-06
+ PS=9.3e-07
mX9/X0/X0/M2 N_X9/X0/7_X9/X0/X0/M2_d N_STATE0_X9/X0/X0/M2_g N_VDD_X9/X0/X0/M2_s
+ N_VDD_X7/X0/X0/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.395e-12 AS=2.79e-12 PD=9.3e-07
+ PS=4.86e-06
mX9/X0/X0/M3 N_VDD_X9/X0/X0/M3_d N_STATE0_X9/X0/X0/M3_g N_X9/X0/7_X9/X0/X0/M3_s
+ N_VDD_X7/X0/X0/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.37e-12 AS=1.395e-12
+ PD=4.58e-06 PS=9.3e-07
mX9/X0/X1/M0 N_X9/8_X9/X0/X1/M0_d N_STATE0_X9/X0/X1/M0_g N_INIT3_X9/X0/X1/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.316e-12 AS=1.288e-12 PD=3.28e-06
+ PS=3.24e-06
mX9/X0/X1/M1 N_X9/8_X9/X0/X1/M1_d N_X9/X0/7_X9/X0/X1/M1_g N_INIT3_X9/X0/X1/M1_s
+ N_VDD_X7/X0/X0/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.88e-12 AS=2.7e-12 PD=4.92e-06
+ PS=4.8e-06
mX9/X0/X2/M0 N_X9/8_X9/X0/X2/M0_d N_X9/X0/7_X9/X0/X2/M0_g N_16_X9/X0/X2/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.316e-12 AS=1.288e-12 PD=3.28e-06
+ PS=3.24e-06
mX9/X0/X2/M1 N_X9/8_X9/X0/X2/M1_d N_STATE0_X9/X0/X2/M1_g N_16_X9/X0/X2/M1_s
+ N_VDD_X7/X0/X0/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.88e-12 AS=2.7e-12 PD=4.92e-06
+ PS=4.8e-06
mX9/X1/X0/M0 N_X9/X1/7_X9/X1/X0/M0_d N_STATE1_X9/X1/X0/M0_g N_VSS_X9/X1/X0/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.1625e-12 AS=2.325e-12 PD=9.3e-07
+ PS=4.36e-06
mX9/X1/X0/M1 N_VSS_X9/X1/X0/M1_d N_STATE1_X9/X1/X0/M1_g N_X9/X1/7_X9/X1/X0/M1_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.95e-12 AS=1.1625e-12 PD=4.06e-06
+ PS=9.3e-07
mX9/X1/X0/M2 N_X9/X1/7_X9/X1/X0/M2_d N_STATE1_X9/X1/X0/M2_g N_VDD_X9/X1/X0/M2_s
+ N_VDD_X7/X0/X0/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.395e-12 AS=2.79e-12 PD=9.3e-07
+ PS=4.86e-06
mX9/X1/X0/M3 N_VDD_X9/X1/X0/M3_d N_STATE1_X9/X1/X0/M3_g N_X9/X1/7_X9/X1/X0/M3_s
+ N_VDD_X7/X0/X0/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.37e-12 AS=1.395e-12
+ PD=4.58e-06 PS=9.3e-07
mX9/X1/X1/M0 N_MO3_X9/X1/X1/M0_d N_STATE1_X9/X1/X1/M0_g N_X9/8_X9/X1/X1/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.316e-12 AS=1.288e-12 PD=3.28e-06
+ PS=3.24e-06
mX9/X1/X1/M1 N_MO3_X9/X1/X1/M1_d N_X9/X1/7_X9/X1/X1/M1_g N_X9/8_X9/X1/X1/M1_s
+ N_VDD_X7/X0/X0/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.88e-12 AS=2.7e-12 PD=4.92e-06
+ PS=4.8e-06
mX9/X1/X2/M0 N_MO3_X9/X1/X2/M0_d N_X9/X1/7_X9/X1/X2/M0_g N_VSS_X9/X1/X2/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.316e-12 AS=1.288e-12 PD=3.28e-06
+ PS=3.24e-06
mX9/X1/X2/M1 N_MO3_X9/X1/X2/M1_d N_STATE1_X9/X1/X2/M1_g N_VSS_X9/X1/X2/M1_s
+ N_VDD_X7/X0/X0/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.88e-12 AS=2.7e-12 PD=4.92e-06
+ PS=4.8e-06
mX10/X0/X0/M0 N_X10/X0/7_X10/X0/X0/M0_d N_STATE0_X10/X0/X0/M0_g
+ N_VSS_X10/X0/X0/M0_s N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.1625e-12
+ AS=2.325e-12 PD=9.3e-07 PS=4.36e-06
mX10/X0/X0/M1 N_VSS_X10/X0/X0/M1_d N_STATE0_X10/X0/X0/M1_g
+ N_X10/X0/7_X10/X0/X0/M1_s N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.95e-12
+ AS=1.1625e-12 PD=4.06e-06 PS=9.3e-07
mX10/X0/X0/M2 N_X10/X0/7_X10/X0/X0/M2_d N_STATE0_X10/X0/X0/M2_g
+ N_VDD_X10/X0/X0/M2_s N_VDD_X2/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.395e-12
+ AS=2.79e-12 PD=9.3e-07 PS=4.86e-06
mX10/X0/X0/M3 N_VDD_X10/X0/X0/M3_d N_STATE0_X10/X0/X0/M3_g
+ N_X10/X0/7_X10/X0/X0/M3_s N_VDD_X2/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.37e-12
+ AS=1.395e-12 PD=4.58e-06 PS=9.3e-07
mX10/X0/X1/M0 N_X10/8_X10/X0/X1/M0_d N_STATE0_X10/X0/X1/M0_g
+ N_INIT1_X10/X0/X1/M0_s N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.316e-12
+ AS=1.288e-12 PD=3.28e-06 PS=3.24e-06
mX10/X0/X1/M1 N_X10/8_X10/X0/X1/M1_d N_X10/X0/7_X10/X0/X1/M1_g
+ N_INIT1_X10/X0/X1/M1_s N_VDD_X2/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.88e-12
+ AS=2.7e-12 PD=4.92e-06 PS=4.8e-06
mX10/X0/X2/M0 N_X10/8_X10/X0/X2/M0_d N_X10/X0/7_X10/X0/X2/M0_g
+ N_10_X10/X0/X2/M0_s N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.316e-12
+ AS=1.288e-12 PD=3.28e-06 PS=3.24e-06
mX10/X0/X2/M1 N_X10/8_X10/X0/X2/M1_d N_STATE0_X10/X0/X2/M1_g N_10_X10/X0/X2/M1_s
+ N_VDD_X2/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.88e-12 AS=2.7e-12 PD=4.92e-06
+ PS=4.8e-06
mX10/X1/X0/M0 N_X10/X1/7_X10/X1/X0/M0_d N_STATE1_X10/X1/X0/M0_g
+ N_VSS_X10/X1/X0/M0_s N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.1625e-12
+ AS=2.325e-12 PD=9.3e-07 PS=4.36e-06
mX10/X1/X0/M1 N_VSS_X10/X1/X0/M1_d N_STATE1_X10/X1/X0/M1_g
+ N_X10/X1/7_X10/X1/X0/M1_s N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.95e-12
+ AS=1.1625e-12 PD=4.06e-06 PS=9.3e-07
mX10/X1/X0/M2 N_X10/X1/7_X10/X1/X0/M2_d N_STATE1_X10/X1/X0/M2_g
+ N_VDD_X10/X1/X0/M2_s N_VDD_X2/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.395e-12
+ AS=2.79e-12 PD=9.3e-07 PS=4.86e-06
mX10/X1/X0/M3 N_VDD_X10/X1/X0/M3_d N_STATE1_X10/X1/X0/M3_g
+ N_X10/X1/7_X10/X1/X0/M3_s N_VDD_X2/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.37e-12
+ AS=1.395e-12 PD=4.58e-06 PS=9.3e-07
mX10/X1/X1/M0 N_MO1_X10/X1/X1/M0_d N_STATE1_X10/X1/X1/M0_g
+ N_X10/8_X10/X1/X1/M0_s N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.316e-12
+ AS=1.288e-12 PD=3.28e-06 PS=3.24e-06
mX10/X1/X1/M1 N_MO1_X10/X1/X1/M1_d N_X10/X1/7_X10/X1/X1/M1_g
+ N_X10/8_X10/X1/X1/M1_s N_VDD_X2/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.88e-12
+ AS=2.7e-12 PD=4.92e-06 PS=4.8e-06
mX10/X1/X2/M0 N_MO1_X10/X1/X2/M0_d N_X10/X1/7_X10/X1/X2/M0_g
+ N_VSS_X10/X1/X2/M0_s N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.316e-12
+ AS=1.288e-12 PD=3.28e-06 PS=3.24e-06
mX10/X1/X2/M1 N_MO1_X10/X1/X2/M1_d N_STATE1_X10/X1/X2/M1_g N_VSS_X10/X1/X2/M1_s
+ N_VDD_X2/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.88e-12 AS=2.7e-12 PD=4.92e-06
+ PS=4.8e-06
mX11/M0 N_X11/6_X11/M0_d N_22_X11/M0_g N_VSS_X11/M0_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=1.036e-12 AS=1.008e-12 PD=2.88e-06 PS=2.84e-06
mX11/M1 N_X11/10_X11/M1_d N_CLK_X11/M1_g N_VSS_X11/M1_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=5.6e-13 AS=9.24e-13 PD=8e-07 PS=2.72e-06
mX11/M2 N_X11/7_X11/M2_d N_X11/6_X11/M2_g N_X11/10_X11/M2_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=1.022e-12 AS=5.6e-13 PD=2.86e-06 PS=8e-07
mX11/M3 N_X11/11_X11/M3_d N_X11/7_X11/M3_g N_VSS_X11/M3_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=5.32e-13 AS=9.8e-13 PD=7.6e-07 PS=2.8e-06
mX11/M4 N_X11/8_X11/M4_d N_CLK_X11/M4_g N_X11/11_X11/M4_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=1.022e-12 AS=5.32e-13 PD=2.86e-06 PS=7.6e-07
mX11/M5 N_X11/9_X11/M5_d N_22_X11/M5_g N_VDD_X11/M5_s N_VDD_X11/X9/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=1.2e-12 AS=2.16e-12 PD=8e-07 PS=4.44e-06
mX11/M6 N_X11/6_X11/M6_d N_CLK_X11/M6_g N_X11/9_X11/M6_s N_VDD_X11/X9/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=2.01e-12 AS=1.2e-12 PD=4.34e-06 PS=8e-07
mX11/M7 N_X11/7_X11/M7_d N_CLK_X11/M7_g N_VDD_X11/M7_s N_VDD_X11/X9/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=2.28e-12 AS=2.1e-12 PD=4.52e-06 PS=4.4e-06
mX11/M8 N_X11/8_X11/M8_d N_X11/7_X11/M8_g N_VDD_X11/M8_s N_VDD_X11/X9/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=2.25e-12 AS=2.13e-12 PD=4.5e-06 PS=4.42e-06
mX11/X9/M0 N_STATE1_X11/X9/M0_d N_X11/8_X11/X9/M0_g N_VSS_X11/X9/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.1625e-12 AS=2.325e-12 PD=9.3e-07
+ PS=4.36e-06
mX11/X9/M1 N_VSS_X11/X9/M1_d N_X11/8_X11/X9/M1_g N_STATE1_X11/X9/M1_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.95e-12 AS=1.1625e-12 PD=4.06e-06
+ PS=9.3e-07
mX11/X9/M2 N_STATE1_X11/X9/M2_d N_X11/8_X11/X9/M2_g N_VDD_X11/X9/M2_s
+ N_VDD_X11/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.395e-12 AS=2.79e-12 PD=9.3e-07
+ PS=4.86e-06
mX11/X9/M3 N_VDD_X11/X9/M3_d N_X11/8_X11/X9/M3_g N_STATE1_X11/X9/M3_s
+ N_VDD_X11/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.37e-12 AS=1.395e-12 PD=4.58e-06
+ PS=9.3e-07
mX12/M0 N_X12/6_X12/M0_d N_23_X12/M0_g N_VSS_X12/M0_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=1.036e-12 AS=1.008e-12 PD=2.88e-06 PS=2.84e-06
mX12/M1 N_X12/10_X12/M1_d N_CLK_X12/M1_g N_VSS_X12/M1_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=5.6e-13 AS=9.24e-13 PD=8e-07 PS=2.72e-06
mX12/M2 N_X12/7_X12/M2_d N_X12/6_X12/M2_g N_X12/10_X12/M2_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=1.022e-12 AS=5.6e-13 PD=2.86e-06 PS=8e-07
mX12/M3 N_X12/11_X12/M3_d N_X12/7_X12/M3_g N_VSS_X12/M3_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=5.32e-13 AS=9.8e-13 PD=7.6e-07 PS=2.8e-06
mX12/M4 N_X12/8_X12/M4_d N_CLK_X12/M4_g N_X12/11_X12/M4_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=1.022e-12 AS=5.32e-13 PD=2.86e-06 PS=7.6e-07
mX12/M5 N_X12/9_X12/M5_d N_23_X12/M5_g N_VDD_X12/M5_s N_VDD_X12/X9/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=1.2e-12 AS=2.16e-12 PD=8e-07 PS=4.44e-06
mX12/M6 N_X12/6_X12/M6_d N_CLK_X12/M6_g N_X12/9_X12/M6_s N_VDD_X12/X9/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=2.01e-12 AS=1.2e-12 PD=4.34e-06 PS=8e-07
mX12/M7 N_X12/7_X12/M7_d N_CLK_X12/M7_g N_VDD_X12/M7_s N_VDD_X12/X9/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=2.28e-12 AS=2.1e-12 PD=4.52e-06 PS=4.4e-06
mX12/M8 N_X12/8_X12/M8_d N_X12/7_X12/M8_g N_VDD_X12/M8_s N_VDD_X12/X9/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=2.25e-12 AS=2.13e-12 PD=4.5e-06 PS=4.42e-06
mX12/X9/M0 N_STATE0_X12/X9/M0_d N_X12/8_X12/X9/M0_g N_VSS_X12/X9/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.1625e-12 AS=2.325e-12 PD=9.3e-07
+ PS=4.36e-06
mX12/X9/M1 N_VSS_X12/X9/M1_d N_X12/8_X12/X9/M1_g N_STATE0_X12/X9/M1_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.95e-12 AS=1.1625e-12 PD=4.06e-06
+ PS=9.3e-07
mX12/X9/M2 N_STATE0_X12/X9/M2_d N_X12/8_X12/X9/M2_g N_VDD_X12/X9/M2_s
+ N_VDD_X12/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.395e-12 AS=2.79e-12 PD=9.3e-07
+ PS=4.86e-06
mX12/X9/M3 N_VDD_X12/X9/M3_d N_X12/8_X12/X9/M3_g N_STATE0_X12/X9/M3_s
+ N_VDD_X12/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.37e-12 AS=1.395e-12 PD=4.58e-06
+ PS=9.3e-07
mX13/X0/M0 N_X13/X0/6_X13/X0/M0_d N_M3_X13/X0/M0_g N_VSS_X13/X0/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.036e-12 AS=1.008e-12 PD=2.88e-06
+ PS=2.84e-06
mX13/X0/M1 N_X13/X0/10_X13/X0/M1_d N_26_X13/X0/M1_g N_VSS_X13/X0/M1_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=5.6e-13 AS=9.24e-13 PD=8e-07
+ PS=2.72e-06
mX13/X0/M2 N_X13/X0/7_X13/X0/M2_d N_X13/X0/6_X13/X0/M2_g N_X13/X0/10_X13/X0/M2_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.022e-12 AS=5.6e-13 PD=2.86e-06
+ PS=8e-07
mX13/X0/M3 N_X13/X0/11_X13/X0/M3_d N_X13/X0/7_X13/X0/M3_g N_VSS_X13/X0/M3_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=5.32e-13 AS=9.8e-13 PD=7.6e-07
+ PS=2.8e-06
mX13/X0/M4 N_X13/X0/8_X13/X0/M4_d N_26_X13/X0/M4_g N_X13/X0/11_X13/X0/M4_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.022e-12 AS=5.32e-13 PD=2.86e-06
+ PS=7.6e-07
mX13/X0/M5 N_X13/X0/9_X13/X0/M5_d N_M3_X13/X0/M5_g N_VDD_X13/X0/M5_s
+ N_VDD_X13/X0/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.2e-12 AS=2.16e-12 PD=8e-07
+ PS=4.44e-06
mX13/X0/M6 N_X13/X0/6_X13/X0/M6_d N_26_X13/X0/M6_g N_X13/X0/9_X13/X0/M6_s
+ N_VDD_X13/X0/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.01e-12 AS=1.2e-12 PD=4.34e-06
+ PS=8e-07
mX13/X0/M7 N_X13/X0/7_X13/X0/M7_d N_26_X13/X0/M7_g N_VDD_X13/X0/M7_s
+ N_VDD_X13/X0/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.28e-12 AS=2.1e-12 PD=4.52e-06
+ PS=4.4e-06
mX13/X0/M8 N_X13/X0/8_X13/X0/M8_d N_X13/X0/7_X13/X0/M8_g N_VDD_X13/X0/M8_s
+ N_VDD_X13/X0/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.25e-12 AS=2.13e-12 PD=4.5e-06
+ PS=4.42e-06
mX13/X0/X9/M0 N_16_X13/X0/X9/M0_d N_X13/X0/8_X13/X0/X9/M0_g N_VSS_X13/X0/X9/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.1625e-12 AS=2.325e-12 PD=9.3e-07
+ PS=4.36e-06
mX13/X0/X9/M1 N_VSS_X13/X0/X9/M1_d N_X13/X0/8_X13/X0/X9/M1_g N_16_X13/X0/X9/M1_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.95e-12 AS=1.1625e-12 PD=4.06e-06
+ PS=9.3e-07
mX13/X0/X9/M2 N_16_X13/X0/X9/M2_d N_X13/X0/8_X13/X0/X9/M2_g N_VDD_X13/X0/X9/M2_s
+ N_VDD_X13/X0/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.395e-12 AS=2.79e-12
+ PD=9.3e-07 PS=4.86e-06
mX13/X0/X9/M3 N_VDD_X13/X0/X9/M3_d N_X13/X0/8_X13/X0/X9/M3_g N_16_X13/X0/X9/M3_s
+ N_VDD_X13/X0/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.37e-12 AS=1.395e-12
+ PD=4.58e-06 PS=9.3e-07
mX13/X1/M0 N_X13/X1/6_X13/X1/M0_d N_M1_X13/X1/M0_g N_VSS_X13/X1/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.036e-12 AS=1.008e-12 PD=2.88e-06
+ PS=2.84e-06
mX13/X1/M1 N_X13/X1/10_X13/X1/M1_d N_26_X13/X1/M1_g N_VSS_X13/X1/M1_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=5.6e-13 AS=9.24e-13 PD=8e-07
+ PS=2.72e-06
mX13/X1/M2 N_X13/X1/7_X13/X1/M2_d N_X13/X1/6_X13/X1/M2_g N_X13/X1/10_X13/X1/M2_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.022e-12 AS=5.6e-13 PD=2.86e-06
+ PS=8e-07
mX13/X1/M3 N_X13/X1/11_X13/X1/M3_d N_X13/X1/7_X13/X1/M3_g N_VSS_X13/X1/M3_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=5.32e-13 AS=9.8e-13 PD=7.6e-07
+ PS=2.8e-06
mX13/X1/M4 N_X13/X1/8_X13/X1/M4_d N_26_X13/X1/M4_g N_X13/X1/11_X13/X1/M4_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.022e-12 AS=5.32e-13 PD=2.86e-06
+ PS=7.6e-07
mX13/X1/M5 N_X13/X1/9_X13/X1/M5_d N_M1_X13/X1/M5_g N_VDD_X13/X1/M5_s
+ N_VDD_X13/X1/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.2e-12 AS=2.16e-12 PD=8e-07
+ PS=4.44e-06
mX13/X1/M6 N_X13/X1/6_X13/X1/M6_d N_26_X13/X1/M6_g N_X13/X1/9_X13/X1/M6_s
+ N_VDD_X13/X1/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.01e-12 AS=1.2e-12 PD=4.34e-06
+ PS=8e-07
mX13/X1/M7 N_X13/X1/7_X13/X1/M7_d N_26_X13/X1/M7_g N_VDD_X13/X1/M7_s
+ N_VDD_X13/X1/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.28e-12 AS=2.1e-12 PD=4.52e-06
+ PS=4.4e-06
mX13/X1/M8 N_X13/X1/8_X13/X1/M8_d N_X13/X1/7_X13/X1/M8_g N_VDD_X13/X1/M8_s
+ N_VDD_X13/X1/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.25e-12 AS=2.13e-12 PD=4.5e-06
+ PS=4.42e-06
mX13/X1/X9/M0 N_10_X13/X1/X9/M0_d N_X13/X1/8_X13/X1/X9/M0_g N_VSS_X13/X1/X9/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.1625e-12 AS=2.325e-12 PD=9.3e-07
+ PS=4.36e-06
mX13/X1/X9/M1 N_VSS_X13/X1/X9/M1_d N_X13/X1/8_X13/X1/X9/M1_g N_10_X13/X1/X9/M1_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.95e-12 AS=1.1625e-12 PD=4.06e-06
+ PS=9.3e-07
mX13/X1/X9/M2 N_10_X13/X1/X9/M2_d N_X13/X1/8_X13/X1/X9/M2_g N_VDD_X13/X1/X9/M2_s
+ N_VDD_X13/X1/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.395e-12 AS=2.79e-12
+ PD=9.3e-07 PS=4.86e-06
mX13/X1/X9/M3 N_VDD_X13/X1/X9/M3_d N_X13/X1/8_X13/X1/X9/M3_g N_10_X13/X1/X9/M3_s
+ N_VDD_X13/X1/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.37e-12 AS=1.395e-12
+ PD=4.58e-06 PS=9.3e-07
mX13/X2/M0 N_X13/X2/6_X13/X2/M0_d N_M2_X13/X2/M0_g N_VSS_X13/X2/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.036e-12 AS=1.008e-12 PD=2.88e-06
+ PS=2.84e-06
mX13/X2/M1 N_X13/X2/10_X13/X2/M1_d N_26_X13/X2/M1_g N_VSS_X13/X2/M1_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=5.6e-13 AS=9.24e-13 PD=8e-07
+ PS=2.72e-06
mX13/X2/M2 N_X13/X2/7_X13/X2/M2_d N_X13/X2/6_X13/X2/M2_g N_X13/X2/10_X13/X2/M2_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.022e-12 AS=5.6e-13 PD=2.86e-06
+ PS=8e-07
mX13/X2/M3 N_X13/X2/11_X13/X2/M3_d N_X13/X2/7_X13/X2/M3_g N_VSS_X13/X2/M3_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=5.32e-13 AS=9.8e-13 PD=7.6e-07
+ PS=2.8e-06
mX13/X2/M4 N_X13/X2/8_X13/X2/M4_d N_26_X13/X2/M4_g N_X13/X2/11_X13/X2/M4_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.022e-12 AS=5.32e-13 PD=2.86e-06
+ PS=7.6e-07
mX13/X2/M5 N_X13/X2/9_X13/X2/M5_d N_M2_X13/X2/M5_g N_VDD_X13/X2/M5_s
+ N_VDD_X13/X2/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.2e-12 AS=2.16e-12 PD=8e-07
+ PS=4.44e-06
mX13/X2/M6 N_X13/X2/6_X13/X2/M6_d N_26_X13/X2/M6_g N_X13/X2/9_X13/X2/M6_s
+ N_VDD_X13/X2/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.01e-12 AS=1.2e-12 PD=4.34e-06
+ PS=8e-07
mX13/X2/M7 N_X13/X2/7_X13/X2/M7_d N_26_X13/X2/M7_g N_VDD_X13/X2/M7_s
+ N_VDD_X13/X2/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.28e-12 AS=2.1e-12 PD=4.52e-06
+ PS=4.4e-06
mX13/X2/M8 N_X13/X2/8_X13/X2/M8_d N_X13/X2/7_X13/X2/M8_g N_VDD_X13/X2/M8_s
+ N_VDD_X13/X2/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.25e-12 AS=2.13e-12 PD=4.5e-06
+ PS=4.42e-06
mX13/X2/X9/M0 N_3_X13/X2/X9/M0_d N_X13/X2/8_X13/X2/X9/M0_g N_VSS_X13/X2/X9/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.1625e-12 AS=2.325e-12 PD=9.3e-07
+ PS=4.36e-06
mX13/X2/X9/M1 N_VSS_X13/X2/X9/M1_d N_X13/X2/8_X13/X2/X9/M1_g N_3_X13/X2/X9/M1_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.95e-12 AS=1.1625e-12 PD=4.06e-06
+ PS=9.3e-07
mX13/X2/X9/M2 N_3_X13/X2/X9/M2_d N_X13/X2/8_X13/X2/X9/M2_g N_VDD_X13/X2/X9/M2_s
+ N_VDD_X13/X2/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.395e-12 AS=2.79e-12
+ PD=9.3e-07 PS=4.86e-06
mX13/X2/X9/M3 N_VDD_X13/X2/X9/M3_d N_X13/X2/8_X13/X2/X9/M3_g N_3_X13/X2/X9/M3_s
+ N_VDD_X13/X2/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.37e-12 AS=1.395e-12
+ PD=4.58e-06 PS=9.3e-07
mX13/X3/M0 N_X13/X3/6_X13/X3/M0_d N_M0_X13/X3/M0_g N_VSS_X13/X3/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.036e-12 AS=1.008e-12 PD=2.88e-06
+ PS=2.84e-06
mX13/X3/M1 N_X13/X3/10_X13/X3/M1_d N_26_X13/X3/M1_g N_VSS_X13/X3/M1_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=5.6e-13 AS=9.24e-13 PD=8e-07
+ PS=2.72e-06
mX13/X3/M2 N_X13/X3/7_X13/X3/M2_d N_X13/X3/6_X13/X3/M2_g N_X13/X3/10_X13/X3/M2_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.022e-12 AS=5.6e-13 PD=2.86e-06
+ PS=8e-07
mX13/X3/M3 N_X13/X3/11_X13/X3/M3_d N_X13/X3/7_X13/X3/M3_g N_VSS_X13/X3/M3_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=5.32e-13 AS=9.8e-13 PD=7.6e-07
+ PS=2.8e-06
mX13/X3/M4 N_X13/X3/8_X13/X3/M4_d N_26_X13/X3/M4_g N_X13/X3/11_X13/X3/M4_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.022e-12 AS=5.32e-13 PD=2.86e-06
+ PS=7.6e-07
mX13/X3/M5 N_X13/X3/9_X13/X3/M5_d N_M0_X13/X3/M5_g N_VDD_X13/X3/M5_s
+ N_VDD_X13/X3/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.2e-12 AS=2.16e-12 PD=8e-07
+ PS=4.44e-06
mX13/X3/M6 N_X13/X3/6_X13/X3/M6_d N_26_X13/X3/M6_g N_X13/X3/9_X13/X3/M6_s
+ N_VDD_X13/X3/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.01e-12 AS=1.2e-12 PD=4.34e-06
+ PS=8e-07
mX13/X3/M7 N_X13/X3/7_X13/X3/M7_d N_26_X13/X3/M7_g N_VDD_X13/X3/M7_s
+ N_VDD_X13/X3/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.28e-12 AS=2.1e-12 PD=4.52e-06
+ PS=4.4e-06
mX13/X3/M8 N_X13/X3/8_X13/X3/M8_d N_X13/X3/7_X13/X3/M8_g N_VDD_X13/X3/M8_s
+ N_VDD_X13/X3/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.25e-12 AS=2.13e-12 PD=4.5e-06
+ PS=4.42e-06
mX13/X3/X9/M0 N_4_X13/X3/X9/M0_d N_X13/X3/8_X13/X3/X9/M0_g N_VSS_X13/X3/X9/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.1625e-12 AS=2.325e-12 PD=9.3e-07
+ PS=4.36e-06
mX13/X3/X9/M1 N_VSS_X13/X3/X9/M1_d N_X13/X3/8_X13/X3/X9/M1_g N_4_X13/X3/X9/M1_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.95e-12 AS=1.1625e-12 PD=4.06e-06
+ PS=9.3e-07
mX13/X3/X9/M2 N_4_X13/X3/X9/M2_d N_X13/X3/8_X13/X3/X9/M2_g N_VDD_X13/X3/X9/M2_s
+ N_VDD_X13/X3/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.395e-12 AS=2.79e-12
+ PD=9.3e-07 PS=4.86e-06
mX13/X3/X9/M3 N_VDD_X13/X3/X9/M3_d N_X13/X3/8_X13/X3/X9/M3_g N_4_X13/X3/X9/M3_s
+ N_VDD_X13/X3/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.37e-12 AS=1.395e-12
+ PD=4.58e-06 PS=9.3e-07
mX14/X0/M0 N_X14/X0/6_X14/X0/M0_d N_14_X14/X0/M0_g N_VSS_X14/X0/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.036e-12 AS=1.008e-12 PD=2.88e-06
+ PS=2.84e-06
mX14/X0/M1 N_X14/X0/10_X14/X0/M1_d N_2_X14/X0/M1_g N_VSS_X14/X0/M1_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=5.6e-13 AS=9.24e-13 PD=8e-07
+ PS=2.72e-06
mX14/X0/M2 N_X14/X0/7_X14/X0/M2_d N_X14/X0/6_X14/X0/M2_g N_X14/X0/10_X14/X0/M2_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.022e-12 AS=5.6e-13 PD=2.86e-06
+ PS=8e-07
mX14/X0/M3 N_X14/X0/11_X14/X0/M3_d N_X14/X0/7_X14/X0/M3_g N_VSS_X14/X0/M3_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=5.32e-13 AS=9.8e-13 PD=7.6e-07
+ PS=2.8e-06
mX14/X0/M4 N_X14/X0/8_X14/X0/M4_d N_2_X14/X0/M4_g N_X14/X0/11_X14/X0/M4_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.022e-12 AS=5.32e-13 PD=2.86e-06
+ PS=7.6e-07
mX14/X0/M5 N_X14/X0/9_X14/X0/M5_d N_14_X14/X0/M5_g N_VDD_X14/X0/M5_s
+ N_VDD_X13/X2/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.2e-12 AS=2.16e-12 PD=8e-07
+ PS=4.44e-06
mX14/X0/M6 N_X14/X0/6_X14/X0/M6_d N_2_X14/X0/M6_g N_X14/X0/9_X14/X0/M6_s
+ N_VDD_X13/X2/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.01e-12 AS=1.2e-12 PD=4.34e-06
+ PS=8e-07
mX14/X0/M7 N_X14/X0/7_X14/X0/M7_d N_2_X14/X0/M7_g N_VDD_X14/X0/M7_s
+ N_VDD_X13/X2/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.28e-12 AS=2.1e-12 PD=4.52e-06
+ PS=4.4e-06
mX14/X0/M8 N_X14/X0/8_X14/X0/M8_d N_X14/X0/7_X14/X0/M8_g N_VDD_X14/X0/M8_s
+ N_VDD_X13/X2/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.25e-12 AS=2.13e-12 PD=4.5e-06
+ PS=4.42e-06
mX14/X0/X9/M0 N_INIT3_X14/X0/X9/M0_d N_X14/X0/8_X14/X0/X9/M0_g
+ N_VSS_X14/X0/X9/M0_s N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.1625e-12
+ AS=2.325e-12 PD=9.3e-07 PS=4.36e-06
mX14/X0/X9/M1 N_VSS_X14/X0/X9/M1_d N_X14/X0/8_X14/X0/X9/M1_g
+ N_INIT3_X14/X0/X9/M1_s N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.95e-12
+ AS=1.1625e-12 PD=4.06e-06 PS=9.3e-07
mX14/X0/X9/M2 N_INIT3_X14/X0/X9/M2_d N_X14/X0/8_X14/X0/X9/M2_g
+ N_VDD_X14/X0/X9/M2_s N_VDD_X13/X2/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.395e-12
+ AS=2.79e-12 PD=9.3e-07 PS=4.86e-06
mX14/X0/X9/M3 N_VDD_X14/X0/X9/M3_d N_X14/X0/8_X14/X0/X9/M3_g
+ N_INIT3_X14/X0/X9/M3_s N_VDD_X13/X2/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.37e-12
+ AS=1.395e-12 PD=4.58e-06 PS=9.3e-07
mX14/X1/M0 N_X14/X1/6_X14/X1/M0_d N_13_X14/X1/M0_g N_VSS_X14/X1/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.036e-12 AS=1.008e-12 PD=2.88e-06
+ PS=2.84e-06
mX14/X1/M1 N_X14/X1/10_X14/X1/M1_d N_2_X14/X1/M1_g N_VSS_X14/X1/M1_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=5.6e-13 AS=9.24e-13 PD=8e-07
+ PS=2.72e-06
mX14/X1/M2 N_X14/X1/7_X14/X1/M2_d N_X14/X1/6_X14/X1/M2_g N_X14/X1/10_X14/X1/M2_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.022e-12 AS=5.6e-13 PD=2.86e-06
+ PS=8e-07
mX14/X1/M3 N_X14/X1/11_X14/X1/M3_d N_X14/X1/7_X14/X1/M3_g N_VSS_X14/X1/M3_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=5.32e-13 AS=9.8e-13 PD=7.6e-07
+ PS=2.8e-06
mX14/X1/M4 N_X14/X1/8_X14/X1/M4_d N_2_X14/X1/M4_g N_X14/X1/11_X14/X1/M4_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.022e-12 AS=5.32e-13 PD=2.86e-06
+ PS=7.6e-07
mX14/X1/M5 N_X14/X1/9_X14/X1/M5_d N_13_X14/X1/M5_g N_VDD_X14/X1/M5_s
+ N_VDD_X13/X3/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.2e-12 AS=2.16e-12 PD=8e-07
+ PS=4.44e-06
mX14/X1/M6 N_X14/X1/6_X14/X1/M6_d N_2_X14/X1/M6_g N_X14/X1/9_X14/X1/M6_s
+ N_VDD_X13/X3/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.01e-12 AS=1.2e-12 PD=4.34e-06
+ PS=8e-07
mX14/X1/M7 N_X14/X1/7_X14/X1/M7_d N_2_X14/X1/M7_g N_VDD_X14/X1/M7_s
+ N_VDD_X13/X3/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.28e-12 AS=2.1e-12 PD=4.52e-06
+ PS=4.4e-06
mX14/X1/M8 N_X14/X1/8_X14/X1/M8_d N_X14/X1/7_X14/X1/M8_g N_VDD_X14/X1/M8_s
+ N_VDD_X13/X3/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.25e-12 AS=2.13e-12 PD=4.5e-06
+ PS=4.42e-06
mX14/X1/X9/M0 N_INIT1_X14/X1/X9/M0_d N_X14/X1/8_X14/X1/X9/M0_g
+ N_VSS_X14/X1/X9/M0_s N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.1625e-12
+ AS=2.325e-12 PD=9.3e-07 PS=4.36e-06
mX14/X1/X9/M1 N_VSS_X14/X1/X9/M1_d N_X14/X1/8_X14/X1/X9/M1_g
+ N_INIT1_X14/X1/X9/M1_s N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.95e-12
+ AS=1.1625e-12 PD=4.06e-06 PS=9.3e-07
mX14/X1/X9/M2 N_INIT1_X14/X1/X9/M2_d N_X14/X1/8_X14/X1/X9/M2_g
+ N_VDD_X14/X1/X9/M2_s N_VDD_X13/X3/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.395e-12
+ AS=2.79e-12 PD=9.3e-07 PS=4.86e-06
mX14/X1/X9/M3 N_VDD_X14/X1/X9/M3_d N_X14/X1/8_X14/X1/X9/M3_g
+ N_INIT1_X14/X1/X9/M3_s N_VDD_X13/X3/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.37e-12
+ AS=1.395e-12 PD=4.58e-06 PS=9.3e-07
mX14/X2/M0 N_X14/X2/6_X14/X2/M0_d N_27_X14/X2/M0_g N_VSS_X14/X2/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.036e-12 AS=1.008e-12 PD=2.88e-06
+ PS=2.84e-06
mX14/X2/M1 N_X14/X2/10_X14/X2/M1_d N_2_X14/X2/M1_g N_VSS_X14/X2/M1_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=5.6e-13 AS=9.24e-13 PD=8e-07
+ PS=2.72e-06
mX14/X2/M2 N_X14/X2/7_X14/X2/M2_d N_X14/X2/6_X14/X2/M2_g N_X14/X2/10_X14/X2/M2_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.022e-12 AS=5.6e-13 PD=2.86e-06
+ PS=8e-07
mX14/X2/M3 N_X14/X2/11_X14/X2/M3_d N_X14/X2/7_X14/X2/M3_g N_VSS_X14/X2/M3_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=5.32e-13 AS=9.8e-13 PD=7.6e-07
+ PS=2.8e-06
mX14/X2/M4 N_X14/X2/8_X14/X2/M4_d N_2_X14/X2/M4_g N_X14/X2/11_X14/X2/M4_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.022e-12 AS=5.32e-13 PD=2.86e-06
+ PS=7.6e-07
mX14/X2/M5 N_X14/X2/9_X14/X2/M5_d N_27_X14/X2/M5_g N_VDD_X14/X2/M5_s
+ N_VDD_X14/X2/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.2e-12 AS=2.16e-12 PD=8e-07
+ PS=4.44e-06
mX14/X2/M6 N_X14/X2/6_X14/X2/M6_d N_2_X14/X2/M6_g N_X14/X2/9_X14/X2/M6_s
+ N_VDD_X14/X2/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.01e-12 AS=1.2e-12 PD=4.34e-06
+ PS=8e-07
mX14/X2/M7 N_X14/X2/7_X14/X2/M7_d N_2_X14/X2/M7_g N_VDD_X14/X2/M7_s
+ N_VDD_X14/X2/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.28e-12 AS=2.1e-12 PD=4.52e-06
+ PS=4.4e-06
mX14/X2/M8 N_X14/X2/8_X14/X2/M8_d N_X14/X2/7_X14/X2/M8_g N_VDD_X14/X2/M8_s
+ N_VDD_X14/X2/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.25e-12 AS=2.13e-12 PD=4.5e-06
+ PS=4.42e-06
mX14/X2/X9/M0 N_INIT2_X14/X2/X9/M0_d N_X14/X2/8_X14/X2/X9/M0_g
+ N_VSS_X14/X2/X9/M0_s N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.1625e-12
+ AS=2.325e-12 PD=9.3e-07 PS=4.36e-06
mX14/X2/X9/M1 N_VSS_X14/X2/X9/M1_d N_X14/X2/8_X14/X2/X9/M1_g
+ N_INIT2_X14/X2/X9/M1_s N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.95e-12
+ AS=1.1625e-12 PD=4.06e-06 PS=9.3e-07
mX14/X2/X9/M2 N_INIT2_X14/X2/X9/M2_d N_X14/X2/8_X14/X2/X9/M2_g
+ N_VDD_X14/X2/X9/M2_s N_VDD_X14/X2/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.395e-12
+ AS=2.79e-12 PD=9.3e-07 PS=4.86e-06
mX14/X2/X9/M3 N_VDD_X14/X2/X9/M3_d N_X14/X2/8_X14/X2/X9/M3_g
+ N_INIT2_X14/X2/X9/M3_s N_VDD_X14/X2/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.37e-12
+ AS=1.395e-12 PD=4.58e-06 PS=9.3e-07
mX14/X3/M0 N_X14/X3/6_X14/X3/M0_d N_5_X14/X3/M0_g N_VSS_X14/X3/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.036e-12 AS=1.008e-12 PD=2.88e-06
+ PS=2.84e-06
mX14/X3/M1 N_X14/X3/10_X14/X3/M1_d N_2_X14/X3/M1_g N_VSS_X14/X3/M1_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=5.6e-13 AS=9.24e-13 PD=8e-07
+ PS=2.72e-06
mX14/X3/M2 N_X14/X3/7_X14/X3/M2_d N_X14/X3/6_X14/X3/M2_g N_X14/X3/10_X14/X3/M2_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.022e-12 AS=5.6e-13 PD=2.86e-06
+ PS=8e-07
mX14/X3/M3 N_X14/X3/11_X14/X3/M3_d N_X14/X3/7_X14/X3/M3_g N_VSS_X14/X3/M3_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=5.32e-13 AS=9.8e-13 PD=7.6e-07
+ PS=2.8e-06
mX14/X3/M4 N_X14/X3/8_X14/X3/M4_d N_2_X14/X3/M4_g N_X14/X3/11_X14/X3/M4_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=1.022e-12 AS=5.32e-13 PD=2.86e-06
+ PS=7.6e-07
mX14/X3/M5 N_X14/X3/9_X14/X3/M5_d N_5_X14/X3/M5_g N_VDD_X14/X3/M5_s
+ N_VDD_X14/X3/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.2e-12 AS=2.16e-12 PD=8e-07
+ PS=4.44e-06
mX14/X3/M6 N_X14/X3/6_X14/X3/M6_d N_2_X14/X3/M6_g N_X14/X3/9_X14/X3/M6_s
+ N_VDD_X14/X3/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.01e-12 AS=1.2e-12 PD=4.34e-06
+ PS=8e-07
mX14/X3/M7 N_X14/X3/7_X14/X3/M7_d N_2_X14/X3/M7_g N_VDD_X14/X3/M7_s
+ N_VDD_X14/X3/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.28e-12 AS=2.1e-12 PD=4.52e-06
+ PS=4.4e-06
mX14/X3/M8 N_X14/X3/8_X14/X3/M8_d N_X14/X3/7_X14/X3/M8_g N_VDD_X14/X3/M8_s
+ N_VDD_X14/X3/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.25e-12 AS=2.13e-12 PD=4.5e-06
+ PS=4.42e-06
mX14/X3/X9/M0 N_INIT0_X14/X3/X9/M0_d N_X14/X3/8_X14/X3/X9/M0_g
+ N_VSS_X14/X3/X9/M0_s N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.1625e-12
+ AS=2.325e-12 PD=9.3e-07 PS=4.36e-06
mX14/X3/X9/M1 N_VSS_X14/X3/X9/M1_d N_X14/X3/8_X14/X3/X9/M1_g
+ N_INIT0_X14/X3/X9/M1_s N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.95e-12
+ AS=1.1625e-12 PD=4.06e-06 PS=9.3e-07
mX14/X3/X9/M2 N_INIT0_X14/X3/X9/M2_d N_X14/X3/8_X14/X3/X9/M2_g
+ N_VDD_X14/X3/X9/M2_s N_VDD_X14/X3/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.395e-12
+ AS=2.79e-12 PD=9.3e-07 PS=4.86e-06
mX14/X3/X9/M3 N_VDD_X14/X3/X9/M3_d N_X14/X3/8_X14/X3/X9/M3_g
+ N_INIT0_X14/X3/X9/M3_s N_VDD_X14/X3/X9/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.37e-12
+ AS=1.395e-12 PD=4.58e-06 PS=9.3e-07
mX15/M0 N_X15/7_X15/M0_d N_STATE1_X15/M0_g N_VSS_X15/M0_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=5.18e-13 AS=1.022e-12 PD=7.4e-07 PS=2.86e-06
mX15/M1 N_X15/6_X15/M1_d N_STATE0_X15/M1_g N_X15/7_X15/M1_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=9.24e-13 AS=5.18e-13 PD=2.72e-06 PS=7.4e-07
mX15/M2 N_X15/6_X15/M2_d N_STATE1_X15/M2_g N_VDD_X15/M2_s N_VDD_X15/X4/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=1.11e-12 AS=2.19e-12 PD=7.4e-07 PS=4.46e-06
mX15/M3 N_VDD_X15/M3_d N_STATE0_X15/M3_g N_X15/6_X15/M3_s N_VDD_X15/X4/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=2.19e-12 AS=1.11e-12 PD=4.46e-06 PS=7.4e-07
mX15/X4/M0 N_2_X15/X4/M0_d N_X15/6_X15/X4/M0_g N_VSS_X15/X4/M0_s N_VSS_X0/M0_b
+ N_18 L=1.8e-07 W=2.5e-06 AD=1.1625e-12 AS=2.325e-12 PD=9.3e-07 PS=4.36e-06
mX15/X4/M1 N_VSS_X15/X4/M1_d N_X15/6_X15/X4/M1_g N_2_X15/X4/M1_s N_VSS_X0/M0_b
+ N_18 L=1.8e-07 W=2.5e-06 AD=1.95e-12 AS=1.1625e-12 PD=4.06e-06 PS=9.3e-07
mX15/X4/M2 N_2_X15/X4/M2_d N_X15/6_X15/X4/M2_g N_VDD_X15/X4/M2_s
+ N_VDD_X15/X4/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.395e-12 AS=2.79e-12 PD=9.3e-07
+ PS=4.86e-06
mX15/X4/M3 N_VDD_X15/X4/M3_d N_X15/6_X15/X4/M3_g N_2_X15/X4/M3_s
+ N_VDD_X15/X4/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.37e-12 AS=1.395e-12 PD=4.58e-06
+ PS=9.3e-07
mX16/M0 N_S3_X16/M0_d N_32_X16/M0_g N_VSS_X16/M0_s N_VSS_X0/M0_b N_18 L=1.8e-07
+ W=1.4e-06 AD=5.18e-13 AS=1.022e-12 PD=7.4e-07 PS=2.86e-06
mX16/M1 N_VSS_X16/M1_d N_24_X16/M1_g N_S3_X16/M1_s N_VSS_X0/M0_b N_18 L=1.8e-07
+ W=1.4e-06 AD=9.24e-13 AS=5.18e-13 PD=2.72e-06 PS=7.4e-07
mX16/M2 N_X16/6_X16/M2_d N_32_X16/M2_g N_VDD_X16/M2_s N_VDD_X16/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=1.11e-12 AS=2.19e-12 PD=7.4e-07 PS=4.46e-06
mX16/M3 N_S3_X16/M3_d N_24_X16/M3_g N_X16/6_X16/M3_s N_VDD_X16/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=2.19e-12 AS=1.11e-12 PD=4.46e-06 PS=7.4e-07
mX17/M0 N_S2_X17/M0_d N_32_X17/M0_g N_VSS_X17/M0_s N_VSS_X0/M0_b N_18 L=1.8e-07
+ W=1.4e-06 AD=5.18e-13 AS=1.022e-12 PD=7.4e-07 PS=2.86e-06
mX17/M1 N_VSS_X17/M1_d N_STATE0_X17/M1_g N_S2_X17/M1_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=9.24e-13 AS=5.18e-13 PD=2.72e-06 PS=7.4e-07
mX17/M2 N_X17/6_X17/M2_d N_32_X17/M2_g N_VDD_X17/M2_s N_VDD_X17/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=1.11e-12 AS=2.19e-12 PD=7.4e-07 PS=4.46e-06
mX17/M3 N_S2_X17/M3_d N_STATE0_X17/M3_g N_X17/6_X17/M3_s N_VDD_X17/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=2.19e-12 AS=1.11e-12 PD=4.46e-06 PS=7.4e-07
mX18/M0 N_S1_X18/M0_d N_STATE1_X18/M0_g N_VSS_X18/M0_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=5.18e-13 AS=1.022e-12 PD=7.4e-07 PS=2.86e-06
mX18/M1 N_VSS_X18/M1_d N_24_X18/M1_g N_S1_X18/M1_s N_VSS_X0/M0_b N_18 L=1.8e-07
+ W=1.4e-06 AD=9.24e-13 AS=5.18e-13 PD=2.72e-06 PS=7.4e-07
mX18/M2 N_X18/6_X18/M2_d N_STATE1_X18/M2_g N_VDD_X18/M2_s N_VDD_X18/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=1.11e-12 AS=2.19e-12 PD=7.4e-07 PS=4.46e-06
mX18/M3 N_S1_X18/M3_d N_24_X18/M3_g N_X18/6_X18/M3_s N_VDD_X18/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=2.19e-12 AS=1.11e-12 PD=4.46e-06 PS=7.4e-07
mX19/M0 N_S0_X19/M0_d N_STATE1_X19/M0_g N_VSS_X19/M0_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=5.18e-13 AS=1.022e-12 PD=7.4e-07 PS=2.86e-06
mX19/M1 N_VSS_X19/M1_d N_STATE0_X19/M1_g N_S0_X19/M1_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=9.24e-13 AS=5.18e-13 PD=2.72e-06 PS=7.4e-07
mX19/M2 N_X19/6_X19/M2_d N_STATE1_X19/M2_g N_VDD_X19/M2_s N_VDD_X19/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=1.11e-12 AS=2.19e-12 PD=7.4e-07 PS=4.46e-06
mX19/M3 N_S0_X19/M3_d N_STATE0_X19/M3_g N_X19/6_X19/M3_s N_VDD_X19/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=2.19e-12 AS=1.11e-12 PD=4.46e-06 PS=7.4e-07
mX20/M0 N_X20/8_X20/M0_d N_33_X20/M0_g N_VSS_X20/M0_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=5.18e-13 AS=1.022e-12 PD=7.4e-07 PS=2.86e-06
mX20/M1 N_X20/9_X20/M1_d N_STATE0_X20/M1_g N_X20/8_X20/M1_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=5.04e-13 AS=5.18e-13 PD=7.2e-07 PS=7.4e-07
mX20/M2 N_X20/7_X20/M2_d N_STORE_X20/M2_g N_X20/9_X20/M2_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=8.4e-13 AS=5.04e-13 PD=2.6e-06 PS=7.2e-07
mX20/M3 N_X20/7_X20/M3_d N_33_X20/M3_g N_VDD_X20/M3_s N_VDD_X20/X6/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=1.11e-12 AS=2.19e-12 PD=7.4e-07 PS=4.46e-06
mX20/M4 N_VDD_X20/M4_d N_STATE0_X20/M4_g N_X20/7_X20/M4_s N_VDD_X20/X6/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=1.08e-12 AS=1.11e-12 PD=7.2e-07 PS=7.4e-07
mX20/M5 N_X20/7_X20/M5_d N_STORE_X20/M5_g N_VDD_X20/M5_s N_VDD_X20/X6/M2_b P_18
+ L=1.8e-07 W=3e-06 AD=2.07e-12 AS=1.08e-12 PD=4.38e-06 PS=7.2e-07
mX20/X6/M0 N_26_X20/X6/M0_d N_X20/7_X20/X6/M0_g N_VSS_X20/X6/M0_s N_VSS_X0/M0_b
+ N_18 L=1.8e-07 W=2.5e-06 AD=1.1625e-12 AS=2.325e-12 PD=9.3e-07 PS=4.36e-06
mX20/X6/M1 N_VSS_X20/X6/M1_d N_X20/7_X20/X6/M1_g N_26_X20/X6/M1_s N_VSS_X0/M0_b
+ N_18 L=1.8e-07 W=2.5e-06 AD=1.95e-12 AS=1.1625e-12 PD=4.06e-06 PS=9.3e-07
mX20/X6/M2 N_26_X20/X6/M2_d N_X20/7_X20/X6/M2_g N_VDD_X20/X6/M2_s
+ N_VDD_X20/X6/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.395e-12 AS=2.79e-12 PD=9.3e-07
+ PS=4.86e-06
mX20/X6/M3 N_VDD_X20/X6/M3_d N_X20/7_X20/X6/M3_g N_26_X20/X6/M3_s
+ N_VDD_X20/X6/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.37e-12 AS=1.395e-12 PD=4.58e-06
+ PS=9.3e-07
mX21/M0 N_X21/23_X21/M0_d N_POWER_X21/M0_g N_VSS_X21/M0_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=5.18e-13 AS=1.022e-12 PD=7.4e-07 PS=2.86e-06
mX21/M1 N_X21/24_X21/M1_d N_X21/16_X21/M1_g N_X21/23_X21/M1_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=5.04e-13 AS=5.18e-13 PD=7.2e-07 PS=7.4e-07
mX21/M2 N_X21/25_X21/M2_d N_STATE0_X21/M2_g N_X21/24_X21/M2_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=5.18e-13 AS=5.04e-13 PD=7.4e-07 PS=7.2e-07
mX21/M3 N_X21/17_X21/M3_d N_STORE_X21/M3_g N_X21/25_X21/M3_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=7.42e-13 AS=5.18e-13 PD=2.46e-06 PS=7.4e-07
mX21/M4 N_X21/20_X21/M4_d N_X21/15_X21/M4_g N_VSS_X21/M4_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=5.18e-13 AS=1.022e-12 PD=7.4e-07 PS=2.86e-06
mX21/M5 N_VSS_X21/M5_d N_X21/14_X21/M5_g N_X21/20_X21/M5_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=5.11e-13 AS=5.18e-13 PD=7.3e-07 PS=7.4e-07
mX21/M6 N_X21/20_X21/M6_d N_X21/10_X21/M6_g N_VSS_X21/M6_s N_VSS_X0/M0_b N_18
+ L=1.8e-07 W=1.4e-06 AD=1.036e-12 AS=5.11e-13 PD=2.88e-06 PS=7.3e-07
mX21/M7 N_X21/17_X21/M7_d N_POWER_X21/M7_g N_VDD_X21/M7_s N_VDD_X21/X18/M2_b
+ P_18 L=1.8e-07 W=3e-06 AD=1.11e-12 AS=2.19e-12 PD=7.4e-07 PS=4.46e-06
mX21/M8 N_VDD_X21/M8_d N_X21/16_X21/M8_g N_X21/17_X21/M8_s N_VDD_X21/X18/M2_b
+ P_18 L=1.8e-07 W=3e-06 AD=1.08e-12 AS=1.11e-12 PD=7.2e-07 PS=7.4e-07
mX21/M9 N_X21/17_X21/M9_d N_STATE0_X21/M9_g N_VDD_X21/M9_s N_VDD_X21/X18/M2_b
+ P_18 L=1.8e-07 W=3e-06 AD=1.11e-12 AS=1.08e-12 PD=7.4e-07 PS=7.2e-07
mX21/M10 N_VDD_X21/M10_d N_STORE_X21/M10_g N_X21/17_X21/M10_s N_VDD_X21/X18/M2_b
+ P_18 L=1.8e-07 W=3e-06 AD=1.8e-12 AS=1.11e-12 PD=4.2e-06 PS=7.4e-07
mX21/M11 N_X21/21_X21/M11_d N_X21/15_X21/M11_g N_VDD_X21/M11_s
+ N_VDD_X21/X20/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.11e-12 AS=2.19e-12 PD=7.4e-07
+ PS=4.46e-06
mX21/M12 N_X21/22_X21/M12_d N_X21/14_X21/M12_g N_X21/21_X21/M12_s
+ N_VDD_X21/X20/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.095e-12 AS=1.11e-12 PD=7.3e-07
+ PS=7.4e-07
mX21/M13 N_X21/20_X21/M13_d N_X21/10_X21/M13_g N_X21/22_X21/M13_s
+ N_VDD_X21/X20/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.19e-12 AS=1.095e-12 PD=4.46e-06
+ PS=7.3e-07
mX21/X14/M0 N_X21/16_X21/X14/M0_d N_STATE1_X21/X14/M0_g N_VSS_X21/X14/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.1625e-12 AS=2.325e-12 PD=9.3e-07
+ PS=4.36e-06
mX21/X14/M1 N_VSS_X21/X14/M1_d N_STATE1_X21/X14/M1_g N_X21/16_X21/X14/M1_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.95e-12 AS=1.1625e-12 PD=4.06e-06
+ PS=9.3e-07
mX21/X14/M2 N_X21/16_X21/X14/M2_d N_STATE1_X21/X14/M2_g N_VDD_X21/X14/M2_s
+ N_VDD_X21/X14/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.395e-12 AS=2.79e-12 PD=9.3e-07
+ PS=4.86e-06
mX21/X14/M3 N_VDD_X21/X14/M3_d N_STATE1_X21/X14/M3_g N_X21/16_X21/X14/M3_s
+ N_VDD_X21/X14/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.37e-12 AS=1.395e-12 PD=4.58e-06
+ PS=9.3e-07
mX21/X15/M0 N_X21/12_X21/X15/M0_d N_STORE_X21/X15/M0_g N_VSS_X21/X15/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.1625e-12 AS=2.325e-12 PD=9.3e-07
+ PS=4.36e-06
mX21/X15/M1 N_VSS_X21/X15/M1_d N_STORE_X21/X15/M1_g N_X21/12_X21/X15/M1_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.95e-12 AS=1.1625e-12 PD=4.06e-06
+ PS=9.3e-07
mX21/X15/M2 N_X21/12_X21/X15/M2_d N_STORE_X21/X15/M2_g N_VDD_X21/X15/M2_s
+ N_VDD_X21/X15/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.395e-12 AS=2.79e-12 PD=9.3e-07
+ PS=4.86e-06
mX21/X15/M3 N_VDD_X21/X15/M3_d N_STORE_X21/X15/M3_g N_X21/12_X21/X15/M3_s
+ N_VDD_X21/X15/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.37e-12 AS=1.395e-12 PD=4.58e-06
+ PS=9.3e-07
mX21/X16/M0 N_X21/9_X21/X16/M0_d N_STATE0_X21/X16/M0_g N_VSS_X21/X16/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.1625e-12 AS=2.325e-12 PD=9.3e-07
+ PS=4.36e-06
mX21/X16/M1 N_VSS_X21/X16/M1_d N_STATE0_X21/X16/M1_g N_X21/9_X21/X16/M1_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.95e-12 AS=1.1625e-12 PD=4.06e-06
+ PS=9.3e-07
mX21/X16/M2 N_X21/9_X21/X16/M2_d N_STATE0_X21/X16/M2_g N_VDD_X21/X16/M2_s
+ N_VDD_X21/X16/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.395e-12 AS=2.79e-12 PD=9.3e-07
+ PS=4.86e-06
mX21/X16/M3 N_VDD_X21/X16/M3_d N_STATE0_X21/X16/M3_g N_X21/9_X21/X16/M3_s
+ N_VDD_X21/X16/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.37e-12 AS=1.395e-12 PD=4.58e-06
+ PS=9.3e-07
mX21/X17/M0 N_X21/11_X21/X17/M0_d N_STATE0_X21/X17/M0_g N_VSS_X21/X17/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.1625e-12 AS=2.325e-12 PD=9.3e-07
+ PS=4.36e-06
mX21/X17/M1 N_VSS_X21/X17/M1_d N_STATE0_X21/X17/M1_g N_X21/11_X21/X17/M1_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.95e-12 AS=1.1625e-12 PD=4.06e-06
+ PS=9.3e-07
mX21/X17/M2 N_X21/11_X21/X17/M2_d N_STATE0_X21/X17/M2_g N_VDD_X21/X17/M2_s
+ N_VDD_X21/X17/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.395e-12 AS=2.79e-12 PD=9.3e-07
+ PS=4.86e-06
mX21/X17/M3 N_VDD_X21/X17/M3_d N_STATE0_X21/X17/M3_g N_X21/11_X21/X17/M3_s
+ N_VDD_X21/X17/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.37e-12 AS=1.395e-12 PD=4.58e-06
+ PS=9.3e-07
mX21/X18/M0 N_X21/13_X21/X18/M0_d N_X21/17_X21/X18/M0_g N_VSS_X21/X18/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.1625e-12 AS=2.325e-12 PD=9.3e-07
+ PS=4.36e-06
mX21/X18/M1 N_VSS_X21/X18/M1_d N_X21/17_X21/X18/M1_g N_X21/13_X21/X18/M1_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.95e-12 AS=1.1625e-12 PD=4.06e-06
+ PS=9.3e-07
mX21/X18/M2 N_X21/13_X21/X18/M2_d N_X21/17_X21/X18/M2_g N_VDD_X21/X18/M2_s
+ N_VDD_X21/X18/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.395e-12 AS=2.79e-12 PD=9.3e-07
+ PS=4.86e-06
mX21/X18/M3 N_VDD_X21/X18/M3_d N_X21/17_X21/X18/M3_g N_X21/13_X21/X18/M3_s
+ N_VDD_X21/X18/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.37e-12 AS=1.395e-12 PD=4.58e-06
+ PS=9.3e-07
mX21/X19/M0 N_22_X21/X19/M0_d N_X21/19_X21/X19/M0_g N_VSS_X21/X19/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.1625e-12 AS=2.325e-12 PD=9.3e-07
+ PS=4.36e-06
mX21/X19/M1 N_VSS_X21/X19/M1_d N_X21/19_X21/X19/M1_g N_22_X21/X19/M1_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.95e-12 AS=1.1625e-12 PD=4.06e-06
+ PS=9.3e-07
mX21/X19/M2 N_22_X21/X19/M2_d N_X21/19_X21/X19/M2_g N_VDD_X21/X19/M2_s
+ N_VDD_X21/X19/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.395e-12 AS=2.79e-12 PD=9.3e-07
+ PS=4.86e-06
mX21/X19/M3 N_VDD_X21/X19/M3_d N_X21/19_X21/X19/M3_g N_22_X21/X19/M3_s
+ N_VDD_X21/X19/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.37e-12 AS=1.395e-12 PD=4.58e-06
+ PS=9.3e-07
mX21/X20/M0 N_23_X21/X20/M0_d N_X21/20_X21/X20/M0_g N_VSS_X21/X20/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.1625e-12 AS=2.325e-12 PD=9.3e-07
+ PS=4.36e-06
mX21/X20/M1 N_VSS_X21/X20/M1_d N_X21/20_X21/X20/M1_g N_23_X21/X20/M1_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.95e-12 AS=1.1625e-12 PD=4.06e-06
+ PS=9.3e-07
mX21/X20/M2 N_23_X21/X20/M2_d N_X21/20_X21/X20/M2_g N_VDD_X21/X20/M2_s
+ N_VDD_X21/X20/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.395e-12 AS=2.79e-12 PD=9.3e-07
+ PS=4.86e-06
mX21/X20/M3 N_VDD_X21/X20/M3_d N_X21/20_X21/X20/M3_g N_23_X21/X20/M3_s
+ N_VDD_X21/X20/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.37e-12 AS=1.395e-12 PD=4.58e-06
+ PS=9.3e-07
mX21/X21/M0 N_X21/X21/7_X21/X21/M0_d N_POWER_X21/X21/M0_g N_VSS_X21/X21/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=5.18e-13 AS=1.022e-12 PD=7.4e-07
+ PS=2.86e-06
mX21/X21/M1 N_X21/X21/6_X21/X21/M1_d N_STATE1_X21/X21/M1_g
+ N_X21/X21/7_X21/X21/M1_s N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=9.24e-13
+ AS=5.18e-13 PD=2.72e-06 PS=7.4e-07
mX21/X21/M2 N_X21/X21/6_X21/X21/M2_d N_POWER_X21/X21/M2_g N_VDD_X21/X21/M2_s
+ N_VDD_X21/X21/X4/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.11e-12 AS=2.19e-12
+ PD=7.4e-07 PS=4.46e-06
mX21/X21/M3 N_VDD_X21/X21/M3_d N_STATE1_X21/X21/M3_g N_X21/X21/6_X21/X21/M3_s
+ N_VDD_X21/X21/X4/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.19e-12 AS=1.11e-12
+ PD=4.46e-06 PS=7.4e-07
mX21/X21/X4/M0 N_X21/15_X21/X21/X4/M0_d N_X21/X21/6_X21/X21/X4/M0_g
+ N_VSS_X21/X21/X4/M0_s N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.1625e-12
+ AS=2.325e-12 PD=9.3e-07 PS=4.36e-06
mX21/X21/X4/M1 N_VSS_X21/X21/X4/M1_d N_X21/X21/6_X21/X21/X4/M1_g
+ N_X21/15_X21/X21/X4/M1_s N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.95e-12
+ AS=1.1625e-12 PD=4.06e-06 PS=9.3e-07
mX21/X21/X4/M2 N_X21/15_X21/X21/X4/M2_d N_X21/X21/6_X21/X21/X4/M2_g
+ N_VDD_X21/X21/X4/M2_s N_VDD_X21/X21/X4/M2_b P_18 L=1.8e-07 W=3e-06
+ AD=1.395e-12 AS=2.79e-12 PD=9.3e-07 PS=4.86e-06
mX21/X21/X4/M3 N_VDD_X21/X21/X4/M3_d N_X21/X21/6_X21/X21/X4/M3_g
+ N_X21/15_X21/X21/X4/M3_s N_VDD_X21/X21/X4/M2_b P_18 L=1.8e-07 W=3e-06
+ AD=2.37e-12 AS=1.395e-12 PD=4.58e-06 PS=9.3e-07
mX21/X22/M0 N_X21/19_X21/X22/M0_d N_X21/18_X21/X22/M0_g N_VSS_X21/X22/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=5.18e-13 AS=1.022e-12 PD=7.4e-07
+ PS=2.86e-06
mX21/X22/M1 N_VSS_X21/X22/M1_d N_X21/13_X21/X22/M1_g N_X21/19_X21/X22/M1_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=9.24e-13 AS=5.18e-13 PD=2.72e-06
+ PS=7.4e-07
mX21/X22/M2 N_X21/X22/6_X21/X22/M2_d N_X21/18_X21/X22/M2_g N_VDD_X21/X22/M2_s
+ N_VDD_X21/X19/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.11e-12 AS=2.19e-12 PD=7.4e-07
+ PS=4.46e-06
mX21/X22/M3 N_X21/19_X21/X22/M3_d N_X21/13_X21/X22/M3_g N_X21/X22/6_X21/X22/M3_s
+ N_VDD_X21/X19/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.19e-12 AS=1.11e-12 PD=4.46e-06
+ PS=7.4e-07
mX21/X23/M0 N_X21/X23/8_X21/X23/M0_d N_POWER_X21/X23/M0_g N_VSS_X21/X23/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=5.18e-13 AS=1.022e-12 PD=7.4e-07
+ PS=2.86e-06
mX21/X23/M1 N_X21/X23/9_X21/X23/M1_d N_STATE1_X21/X23/M1_g
+ N_X21/X23/8_X21/X23/M1_s N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=5.04e-13
+ AS=5.18e-13 PD=7.2e-07 PS=7.4e-07
mX21/X23/M2 N_X21/X23/7_X21/X23/M2_d N_X21/9_X21/X23/M2_g
+ N_X21/X23/9_X21/X23/M2_s N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=8.4e-13
+ AS=5.04e-13 PD=2.6e-06 PS=7.2e-07
mX21/X23/M3 N_X21/X23/7_X21/X23/M3_d N_POWER_X21/X23/M3_g N_VDD_X21/X23/M3_s
+ N_VDD_X21/X19/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.11e-12 AS=2.19e-12 PD=7.4e-07
+ PS=4.46e-06
mX21/X23/M4 N_VDD_X21/X23/M4_d N_STATE1_X21/X23/M4_g N_X21/X23/7_X21/X23/M4_s
+ N_VDD_X21/X19/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.08e-12 AS=1.11e-12 PD=7.2e-07
+ PS=7.4e-07
mX21/X23/M5 N_X21/X23/7_X21/X23/M5_d N_X21/9_X21/X23/M5_g N_VDD_X21/X23/M5_s
+ N_VDD_X21/X19/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.07e-12 AS=1.08e-12 PD=4.38e-06
+ PS=7.2e-07
mX21/X23/X6/M0 N_X21/18_X21/X23/X6/M0_d N_X21/X23/7_X21/X23/X6/M0_g
+ N_VSS_X21/X23/X6/M0_s N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.1625e-12
+ AS=2.325e-12 PD=9.3e-07 PS=4.36e-06
mX21/X23/X6/M1 N_VSS_X21/X23/X6/M1_d N_X21/X23/7_X21/X23/X6/M1_g
+ N_X21/18_X21/X23/X6/M1_s N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.95e-12
+ AS=1.1625e-12 PD=4.06e-06 PS=9.3e-07
mX21/X23/X6/M2 N_X21/18_X21/X23/X6/M2_d N_X21/X23/7_X21/X23/X6/M2_g
+ N_VDD_X21/X23/X6/M2_s N_VDD_X21/X19/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.395e-12
+ AS=2.79e-12 PD=9.3e-07 PS=4.86e-06
mX21/X23/X6/M3 N_VDD_X21/X23/X6/M3_d N_X21/X23/7_X21/X23/X6/M3_g
+ N_X21/18_X21/X23/X6/M3_s N_VDD_X21/X19/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.37e-12
+ AS=1.395e-12 PD=4.58e-06 PS=9.3e-07
mX21/X24/M0 N_X21/X24/8_X21/X24/M0_d N_POWER_X21/X24/M0_g N_VSS_X21/X24/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=5.18e-13 AS=1.022e-12 PD=7.4e-07
+ PS=2.86e-06
mX21/X24/M1 N_X21/X24/9_X21/X24/M1_d N_X21/11_X21/X24/M1_g
+ N_X21/X24/8_X21/X24/M1_s N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=5.04e-13
+ AS=5.18e-13 PD=7.2e-07 PS=7.4e-07
mX21/X24/M2 N_X21/X24/7_X21/X24/M2_d N_STORE_X21/X24/M2_g
+ N_X21/X24/9_X21/X24/M2_s N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=8.4e-13
+ AS=5.04e-13 PD=2.6e-06 PS=7.2e-07
mX21/X24/M3 N_X21/X24/7_X21/X24/M3_d N_POWER_X21/X24/M3_g N_VDD_X21/X24/M3_s
+ N_VDD_X21/X20/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.11e-12 AS=2.19e-12 PD=7.4e-07
+ PS=4.46e-06
mX21/X24/M4 N_VDD_X21/X24/M4_d N_X21/11_X21/X24/M4_g N_X21/X24/7_X21/X24/M4_s
+ N_VDD_X21/X20/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.08e-12 AS=1.11e-12 PD=7.2e-07
+ PS=7.4e-07
mX21/X24/M5 N_X21/X24/7_X21/X24/M5_d N_STORE_X21/X24/M5_g N_VDD_X21/X24/M5_s
+ N_VDD_X21/X20/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.07e-12 AS=1.08e-12 PD=4.38e-06
+ PS=7.2e-07
mX21/X24/X6/M0 N_X21/14_X21/X24/X6/M0_d N_X21/X24/7_X21/X24/X6/M0_g
+ N_VSS_X21/X24/X6/M0_s N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.1625e-12
+ AS=2.325e-12 PD=9.3e-07 PS=4.36e-06
mX21/X24/X6/M1 N_VSS_X21/X24/X6/M1_d N_X21/X24/7_X21/X24/X6/M1_g
+ N_X21/14_X21/X24/X6/M1_s N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.95e-12
+ AS=1.1625e-12 PD=4.06e-06 PS=9.3e-07
mX21/X24/X6/M2 N_X21/14_X21/X24/X6/M2_d N_X21/X24/7_X21/X24/X6/M2_g
+ N_VDD_X21/X24/X6/M2_s N_VDD_X21/X20/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.395e-12
+ AS=2.79e-12 PD=9.3e-07 PS=4.86e-06
mX21/X24/X6/M3 N_VDD_X21/X24/X6/M3_d N_X21/X24/7_X21/X24/X6/M3_g
+ N_X21/14_X21/X24/X6/M3_s N_VDD_X21/X20/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.37e-12
+ AS=1.395e-12 PD=4.58e-06 PS=9.3e-07
mX21/X25/M0 N_X21/X25/8_X21/X25/M0_d N_POWER_X21/X25/M0_g N_VSS_X21/X25/M0_s
+ N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=5.18e-13 AS=1.022e-12 PD=7.4e-07
+ PS=2.86e-06
mX21/X25/M1 N_X21/X25/9_X21/X25/M1_d N_STATE0_X21/X25/M1_g
+ N_X21/X25/8_X21/X25/M1_s N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=5.04e-13
+ AS=5.18e-13 PD=7.2e-07 PS=7.4e-07
mX21/X25/M2 N_X21/X25/7_X21/X25/M2_d N_X21/12_X21/X25/M2_g
+ N_X21/X25/9_X21/X25/M2_s N_VSS_X0/M0_b N_18 L=1.8e-07 W=1.4e-06 AD=8.4e-13
+ AS=5.04e-13 PD=2.6e-06 PS=7.2e-07
mX21/X25/M3 N_X21/X25/7_X21/X25/M3_d N_POWER_X21/X25/M3_g N_VDD_X21/X25/M3_s
+ N_VDD_X21/X21/X4/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.11e-12 AS=2.19e-12
+ PD=7.4e-07 PS=4.46e-06
mX21/X25/M4 N_VDD_X21/X25/M4_d N_STATE0_X21/X25/M4_g N_X21/X25/7_X21/X25/M4_s
+ N_VDD_X21/X21/X4/M2_b P_18 L=1.8e-07 W=3e-06 AD=1.08e-12 AS=1.11e-12
+ PD=7.2e-07 PS=7.4e-07
mX21/X25/M5 N_X21/X25/7_X21/X25/M5_d N_X21/12_X21/X25/M5_g N_VDD_X21/X25/M5_s
+ N_VDD_X21/X21/X4/M2_b P_18 L=1.8e-07 W=3e-06 AD=2.07e-12 AS=1.08e-12
+ PD=4.38e-06 PS=7.2e-07
mX21/X25/X6/M0 N_X21/10_X21/X25/X6/M0_d N_X21/X25/7_X21/X25/X6/M0_g
+ N_VSS_X21/X25/X6/M0_s N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.1625e-12
+ AS=2.325e-12 PD=9.3e-07 PS=4.36e-06
mX21/X25/X6/M1 N_VSS_X21/X25/X6/M1_d N_X21/X25/7_X21/X25/X6/M1_g
+ N_X21/10_X21/X25/X6/M1_s N_VSS_X0/M0_b N_18 L=1.8e-07 W=2.5e-06 AD=1.95e-12
+ AS=1.1625e-12 PD=4.06e-06 PS=9.3e-07
mX21/X25/X6/M2 N_X21/10_X21/X25/X6/M2_d N_X21/X25/7_X21/X25/X6/M2_g
+ N_VDD_X21/X25/X6/M2_s N_VDD_X21/X21/X4/M2_b P_18 L=1.8e-07 W=3e-06
+ AD=1.395e-12 AS=2.79e-12 PD=9.3e-07 PS=4.86e-06
mX21/X25/X6/M3 N_VDD_X21/X25/X6/M3_d N_X21/X25/7_X21/X25/X6/M3_g
+ N_X21/10_X21/X25/X6/M3_s N_VDD_X21/X21/X4/M2_b P_18 L=1.8e-07 W=3e-06
+ AD=2.37e-12 AS=1.395e-12 PD=4.58e-06 PS=9.3e-07
*
.include "Coin_bank.pex.sp.COIN_BANK.pxi"
*
.ends
*
*
